
module InstBufRename ( reset, clk, flush_i, stall_i, instBufferReady_i, 
        decodedPacket0_i, decodedPacket1_i, decodedPacket2_i, decodedPacket3_i, 
        branchCount_i, instBufferReady_o, decodedPacket0_o, decodedPacket1_o, 
        decodedPacket2_o, decodedPacket3_o, branchCount_o );
  input [125:0] decodedPacket0_i;
  input [125:0] decodedPacket1_i;
  input [125:0] decodedPacket2_i;
  input [125:0] decodedPacket3_i;
  input [2:0] branchCount_i;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  output [125:0] decodedPacket2_o;
  output [125:0] decodedPacket3_o;
  output [2:0] branchCount_o;
  input reset, clk, flush_i, stall_i, instBufferReady_i;
  output instBufferReady_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  DFFX1 \branchCount_o_reg[2]  ( .D(n510), .CLK(clk), .Q(branchCount_o[2]) );
  DFFX1 \branchCount_o_reg[1]  ( .D(n509), .CLK(clk), .Q(branchCount_o[1]) );
  DFFX1 \branchCount_o_reg[0]  ( .D(n508), .CLK(clk), .Q(branchCount_o[0]) );
  DFFX1 instBufferReady_o_reg ( .D(n507), .CLK(clk), .Q(instBufferReady_o) );
  DFFX1 \decodedPacket0_o_reg[125]  ( .D(n506), .CLK(clk), .Q(
        decodedPacket0_o[125]) );
  DFFX1 \decodedPacket0_o_reg[124]  ( .D(n505), .CLK(clk), .Q(
        decodedPacket0_o[124]) );
  DFFX1 \decodedPacket0_o_reg[123]  ( .D(n504), .CLK(clk), .Q(
        decodedPacket0_o[123]) );
  DFFX1 \decodedPacket0_o_reg[122]  ( .D(n503), .CLK(clk), .Q(
        decodedPacket0_o[122]) );
  DFFX1 \decodedPacket0_o_reg[121]  ( .D(n502), .CLK(clk), .Q(
        decodedPacket0_o[121]) );
  DFFX1 \decodedPacket0_o_reg[120]  ( .D(n501), .CLK(clk), .Q(
        decodedPacket0_o[120]) );
  DFFX1 \decodedPacket0_o_reg[119]  ( .D(n500), .CLK(clk), .Q(
        decodedPacket0_o[119]) );
  DFFX1 \decodedPacket0_o_reg[118]  ( .D(n499), .CLK(clk), .Q(
        decodedPacket0_o[118]) );
  DFFX1 \decodedPacket0_o_reg[117]  ( .D(n498), .CLK(clk), .Q(
        decodedPacket0_o[117]) );
  DFFX1 \decodedPacket0_o_reg[116]  ( .D(n497), .CLK(clk), .Q(
        decodedPacket0_o[116]) );
  DFFX1 \decodedPacket0_o_reg[115]  ( .D(n496), .CLK(clk), .Q(
        decodedPacket0_o[115]) );
  DFFX1 \decodedPacket0_o_reg[114]  ( .D(n495), .CLK(clk), .Q(
        decodedPacket0_o[114]) );
  DFFX1 \decodedPacket0_o_reg[113]  ( .D(n494), .CLK(clk), .Q(
        decodedPacket0_o[113]) );
  DFFX1 \decodedPacket0_o_reg[112]  ( .D(n493), .CLK(clk), .Q(
        decodedPacket0_o[112]) );
  DFFX1 \decodedPacket0_o_reg[111]  ( .D(n492), .CLK(clk), .Q(
        decodedPacket0_o[111]) );
  DFFX1 \decodedPacket0_o_reg[110]  ( .D(n491), .CLK(clk), .Q(
        decodedPacket0_o[110]) );
  DFFX1 \decodedPacket0_o_reg[109]  ( .D(n490), .CLK(clk), .Q(
        decodedPacket0_o[109]) );
  DFFX1 \decodedPacket0_o_reg[108]  ( .D(n489), .CLK(clk), .Q(
        decodedPacket0_o[108]) );
  DFFX1 \decodedPacket0_o_reg[107]  ( .D(n488), .CLK(clk), .Q(
        decodedPacket0_o[107]) );
  DFFX1 \decodedPacket0_o_reg[106]  ( .D(n487), .CLK(clk), .Q(
        decodedPacket0_o[106]) );
  DFFX1 \decodedPacket0_o_reg[105]  ( .D(n486), .CLK(clk), .Q(
        decodedPacket0_o[105]) );
  DFFX1 \decodedPacket0_o_reg[104]  ( .D(n485), .CLK(clk), .Q(
        decodedPacket0_o[104]) );
  DFFX1 \decodedPacket0_o_reg[103]  ( .D(n484), .CLK(clk), .Q(
        decodedPacket0_o[103]) );
  DFFX1 \decodedPacket0_o_reg[102]  ( .D(n483), .CLK(clk), .Q(
        decodedPacket0_o[102]) );
  DFFX1 \decodedPacket0_o_reg[101]  ( .D(n482), .CLK(clk), .Q(
        decodedPacket0_o[101]) );
  DFFX1 \decodedPacket0_o_reg[100]  ( .D(n481), .CLK(clk), .Q(
        decodedPacket0_o[100]) );
  DFFX1 \decodedPacket0_o_reg[99]  ( .D(n480), .CLK(clk), .Q(
        decodedPacket0_o[99]) );
  DFFX1 \decodedPacket0_o_reg[98]  ( .D(n479), .CLK(clk), .Q(
        decodedPacket0_o[98]) );
  DFFX1 \decodedPacket0_o_reg[97]  ( .D(n478), .CLK(clk), .Q(
        decodedPacket0_o[97]) );
  DFFX1 \decodedPacket0_o_reg[96]  ( .D(n477), .CLK(clk), .Q(
        decodedPacket0_o[96]) );
  DFFX1 \decodedPacket0_o_reg[95]  ( .D(n476), .CLK(clk), .Q(
        decodedPacket0_o[95]) );
  DFFX1 \decodedPacket0_o_reg[94]  ( .D(n475), .CLK(clk), .Q(
        decodedPacket0_o[94]) );
  DFFX1 \decodedPacket0_o_reg[93]  ( .D(n474), .CLK(clk), .Q(
        decodedPacket0_o[93]) );
  DFFX1 \decodedPacket0_o_reg[92]  ( .D(n473), .CLK(clk), .Q(
        decodedPacket0_o[92]) );
  DFFX1 \decodedPacket0_o_reg[91]  ( .D(n472), .CLK(clk), .Q(
        decodedPacket0_o[91]) );
  DFFX1 \decodedPacket0_o_reg[90]  ( .D(n471), .CLK(clk), .Q(
        decodedPacket0_o[90]) );
  DFFX1 \decodedPacket0_o_reg[89]  ( .D(n470), .CLK(clk), .Q(
        decodedPacket0_o[89]) );
  DFFX1 \decodedPacket0_o_reg[88]  ( .D(n469), .CLK(clk), .Q(
        decodedPacket0_o[88]) );
  DFFX1 \decodedPacket0_o_reg[87]  ( .D(n468), .CLK(clk), .Q(
        decodedPacket0_o[87]) );
  DFFX1 \decodedPacket0_o_reg[86]  ( .D(n467), .CLK(clk), .Q(
        decodedPacket0_o[86]) );
  DFFX1 \decodedPacket0_o_reg[85]  ( .D(n466), .CLK(clk), .Q(
        decodedPacket0_o[85]) );
  DFFX1 \decodedPacket0_o_reg[84]  ( .D(n465), .CLK(clk), .Q(
        decodedPacket0_o[84]) );
  DFFX1 \decodedPacket0_o_reg[83]  ( .D(n464), .CLK(clk), .Q(
        decodedPacket0_o[83]) );
  DFFX1 \decodedPacket0_o_reg[82]  ( .D(n463), .CLK(clk), .Q(
        decodedPacket0_o[82]) );
  DFFX1 \decodedPacket0_o_reg[81]  ( .D(n462), .CLK(clk), .Q(
        decodedPacket0_o[81]) );
  DFFX1 \decodedPacket0_o_reg[80]  ( .D(n461), .CLK(clk), .Q(
        decodedPacket0_o[80]) );
  DFFX1 \decodedPacket0_o_reg[79]  ( .D(n460), .CLK(clk), .Q(
        decodedPacket0_o[79]) );
  DFFX1 \decodedPacket0_o_reg[78]  ( .D(n459), .CLK(clk), .Q(
        decodedPacket0_o[78]) );
  DFFX1 \decodedPacket0_o_reg[77]  ( .D(n458), .CLK(clk), .Q(
        decodedPacket0_o[77]) );
  DFFX1 \decodedPacket0_o_reg[76]  ( .D(n457), .CLK(clk), .Q(
        decodedPacket0_o[76]) );
  DFFX1 \decodedPacket0_o_reg[75]  ( .D(n456), .CLK(clk), .Q(
        decodedPacket0_o[75]) );
  DFFX1 \decodedPacket0_o_reg[74]  ( .D(n455), .CLK(clk), .Q(
        decodedPacket0_o[74]) );
  DFFX1 \decodedPacket0_o_reg[73]  ( .D(n454), .CLK(clk), .Q(
        decodedPacket0_o[73]) );
  DFFX1 \decodedPacket0_o_reg[72]  ( .D(n453), .CLK(clk), .Q(
        decodedPacket0_o[72]) );
  DFFX1 \decodedPacket0_o_reg[71]  ( .D(n452), .CLK(clk), .Q(
        decodedPacket0_o[71]) );
  DFFX1 \decodedPacket0_o_reg[70]  ( .D(n451), .CLK(clk), .Q(
        decodedPacket0_o[70]) );
  DFFX1 \decodedPacket0_o_reg[69]  ( .D(n450), .CLK(clk), .Q(
        decodedPacket0_o[69]) );
  DFFX1 \decodedPacket0_o_reg[68]  ( .D(n449), .CLK(clk), .Q(
        decodedPacket0_o[68]) );
  DFFX1 \decodedPacket0_o_reg[67]  ( .D(n448), .CLK(clk), .Q(
        decodedPacket0_o[67]) );
  DFFX1 \decodedPacket0_o_reg[66]  ( .D(n447), .CLK(clk), .Q(
        decodedPacket0_o[66]) );
  DFFX1 \decodedPacket0_o_reg[65]  ( .D(n446), .CLK(clk), .Q(
        decodedPacket0_o[65]) );
  DFFX1 \decodedPacket0_o_reg[64]  ( .D(n445), .CLK(clk), .Q(
        decodedPacket0_o[64]) );
  DFFX1 \decodedPacket0_o_reg[63]  ( .D(n444), .CLK(clk), .Q(
        decodedPacket0_o[63]) );
  DFFX1 \decodedPacket0_o_reg[62]  ( .D(n443), .CLK(clk), .Q(
        decodedPacket0_o[62]) );
  DFFX1 \decodedPacket0_o_reg[61]  ( .D(n442), .CLK(clk), .Q(
        decodedPacket0_o[61]) );
  DFFX1 \decodedPacket0_o_reg[60]  ( .D(n441), .CLK(clk), .Q(
        decodedPacket0_o[60]) );
  DFFX1 \decodedPacket0_o_reg[59]  ( .D(n440), .CLK(clk), .Q(
        decodedPacket0_o[59]) );
  DFFX1 \decodedPacket0_o_reg[58]  ( .D(n439), .CLK(clk), .Q(
        decodedPacket0_o[58]) );
  DFFX1 \decodedPacket0_o_reg[57]  ( .D(n438), .CLK(clk), .Q(
        decodedPacket0_o[57]) );
  DFFX1 \decodedPacket0_o_reg[56]  ( .D(n437), .CLK(clk), .Q(
        decodedPacket0_o[56]) );
  DFFX1 \decodedPacket0_o_reg[55]  ( .D(n436), .CLK(clk), .Q(
        decodedPacket0_o[55]) );
  DFFX1 \decodedPacket0_o_reg[54]  ( .D(n435), .CLK(clk), .Q(
        decodedPacket0_o[54]) );
  DFFX1 \decodedPacket0_o_reg[53]  ( .D(n434), .CLK(clk), .Q(
        decodedPacket0_o[53]) );
  DFFX1 \decodedPacket0_o_reg[52]  ( .D(n433), .CLK(clk), .Q(
        decodedPacket0_o[52]) );
  DFFX1 \decodedPacket0_o_reg[51]  ( .D(n432), .CLK(clk), .Q(
        decodedPacket0_o[51]) );
  DFFX1 \decodedPacket0_o_reg[50]  ( .D(n431), .CLK(clk), .Q(
        decodedPacket0_o[50]) );
  DFFX1 \decodedPacket0_o_reg[49]  ( .D(n430), .CLK(clk), .Q(
        decodedPacket0_o[49]) );
  DFFX1 \decodedPacket0_o_reg[48]  ( .D(n429), .CLK(clk), .Q(
        decodedPacket0_o[48]) );
  DFFX1 \decodedPacket0_o_reg[47]  ( .D(n428), .CLK(clk), .Q(
        decodedPacket0_o[47]) );
  DFFX1 \decodedPacket0_o_reg[46]  ( .D(n427), .CLK(clk), .Q(
        decodedPacket0_o[46]) );
  DFFX1 \decodedPacket0_o_reg[45]  ( .D(n426), .CLK(clk), .Q(
        decodedPacket0_o[45]) );
  DFFX1 \decodedPacket0_o_reg[44]  ( .D(n425), .CLK(clk), .Q(
        decodedPacket0_o[44]) );
  DFFX1 \decodedPacket0_o_reg[43]  ( .D(n424), .CLK(clk), .Q(
        decodedPacket0_o[43]) );
  DFFX1 \decodedPacket0_o_reg[42]  ( .D(n423), .CLK(clk), .Q(
        decodedPacket0_o[42]) );
  DFFX1 \decodedPacket0_o_reg[41]  ( .D(n422), .CLK(clk), .Q(
        decodedPacket0_o[41]) );
  DFFX1 \decodedPacket0_o_reg[40]  ( .D(n421), .CLK(clk), .Q(
        decodedPacket0_o[40]) );
  DFFX1 \decodedPacket0_o_reg[39]  ( .D(n420), .CLK(clk), .Q(
        decodedPacket0_o[39]) );
  DFFX1 \decodedPacket0_o_reg[38]  ( .D(n419), .CLK(clk), .Q(
        decodedPacket0_o[38]) );
  DFFX1 \decodedPacket0_o_reg[37]  ( .D(n418), .CLK(clk), .Q(
        decodedPacket0_o[37]) );
  DFFX1 \decodedPacket0_o_reg[36]  ( .D(n417), .CLK(clk), .Q(
        decodedPacket0_o[36]) );
  DFFX1 \decodedPacket0_o_reg[35]  ( .D(n416), .CLK(clk), .Q(
        decodedPacket0_o[35]) );
  DFFX1 \decodedPacket0_o_reg[34]  ( .D(n415), .CLK(clk), .Q(
        decodedPacket0_o[34]) );
  DFFX1 \decodedPacket0_o_reg[33]  ( .D(n414), .CLK(clk), .Q(
        decodedPacket0_o[33]) );
  DFFX1 \decodedPacket0_o_reg[32]  ( .D(n413), .CLK(clk), .Q(
        decodedPacket0_o[32]) );
  DFFX1 \decodedPacket0_o_reg[31]  ( .D(n412), .CLK(clk), .Q(
        decodedPacket0_o[31]) );
  DFFX1 \decodedPacket0_o_reg[30]  ( .D(n411), .CLK(clk), .Q(
        decodedPacket0_o[30]) );
  DFFX1 \decodedPacket0_o_reg[29]  ( .D(n410), .CLK(clk), .Q(
        decodedPacket0_o[29]) );
  DFFX1 \decodedPacket0_o_reg[28]  ( .D(n409), .CLK(clk), .Q(
        decodedPacket0_o[28]) );
  DFFX1 \decodedPacket0_o_reg[27]  ( .D(n408), .CLK(clk), .Q(
        decodedPacket0_o[27]) );
  DFFX1 \decodedPacket0_o_reg[26]  ( .D(n407), .CLK(clk), .Q(
        decodedPacket0_o[26]) );
  DFFX1 \decodedPacket0_o_reg[25]  ( .D(n406), .CLK(clk), .Q(
        decodedPacket0_o[25]) );
  DFFX1 \decodedPacket0_o_reg[24]  ( .D(n405), .CLK(clk), .Q(
        decodedPacket0_o[24]) );
  DFFX1 \decodedPacket0_o_reg[23]  ( .D(n404), .CLK(clk), .Q(
        decodedPacket0_o[23]) );
  DFFX1 \decodedPacket0_o_reg[22]  ( .D(n403), .CLK(clk), .Q(
        decodedPacket0_o[22]) );
  DFFX1 \decodedPacket0_o_reg[21]  ( .D(n402), .CLK(clk), .Q(
        decodedPacket0_o[21]) );
  DFFX1 \decodedPacket0_o_reg[20]  ( .D(n401), .CLK(clk), .Q(
        decodedPacket0_o[20]) );
  DFFX1 \decodedPacket0_o_reg[19]  ( .D(n400), .CLK(clk), .Q(
        decodedPacket0_o[19]) );
  DFFX1 \decodedPacket0_o_reg[18]  ( .D(n399), .CLK(clk), .Q(
        decodedPacket0_o[18]) );
  DFFX1 \decodedPacket0_o_reg[17]  ( .D(n398), .CLK(clk), .Q(
        decodedPacket0_o[17]) );
  DFFX1 \decodedPacket0_o_reg[16]  ( .D(n397), .CLK(clk), .Q(
        decodedPacket0_o[16]) );
  DFFX1 \decodedPacket0_o_reg[15]  ( .D(n396), .CLK(clk), .Q(
        decodedPacket0_o[15]) );
  DFFX1 \decodedPacket0_o_reg[14]  ( .D(n395), .CLK(clk), .Q(
        decodedPacket0_o[14]) );
  DFFX1 \decodedPacket0_o_reg[13]  ( .D(n394), .CLK(clk), .Q(
        decodedPacket0_o[13]) );
  DFFX1 \decodedPacket0_o_reg[12]  ( .D(n393), .CLK(clk), .Q(
        decodedPacket0_o[12]) );
  DFFX1 \decodedPacket0_o_reg[11]  ( .D(n392), .CLK(clk), .Q(
        decodedPacket0_o[11]) );
  DFFX1 \decodedPacket0_o_reg[10]  ( .D(n391), .CLK(clk), .Q(
        decodedPacket0_o[10]) );
  DFFX1 \decodedPacket0_o_reg[9]  ( .D(n390), .CLK(clk), .Q(
        decodedPacket0_o[9]) );
  DFFX1 \decodedPacket0_o_reg[8]  ( .D(n389), .CLK(clk), .Q(
        decodedPacket0_o[8]) );
  DFFX1 \decodedPacket0_o_reg[7]  ( .D(n388), .CLK(clk), .Q(
        decodedPacket0_o[7]) );
  DFFX1 \decodedPacket0_o_reg[6]  ( .D(n387), .CLK(clk), .Q(
        decodedPacket0_o[6]) );
  DFFX1 \decodedPacket0_o_reg[5]  ( .D(n386), .CLK(clk), .Q(
        decodedPacket0_o[5]) );
  DFFX1 \decodedPacket0_o_reg[4]  ( .D(n385), .CLK(clk), .Q(
        decodedPacket0_o[4]) );
  DFFX1 \decodedPacket0_o_reg[3]  ( .D(n384), .CLK(clk), .Q(
        decodedPacket0_o[3]) );
  DFFX1 \decodedPacket0_o_reg[2]  ( .D(n383), .CLK(clk), .Q(
        decodedPacket0_o[2]) );
  DFFX1 \decodedPacket0_o_reg[1]  ( .D(n382), .CLK(clk), .Q(
        decodedPacket0_o[1]) );
  DFFX1 \decodedPacket0_o_reg[0]  ( .D(n381), .CLK(clk), .Q(
        decodedPacket0_o[0]) );
  DFFX1 \decodedPacket1_o_reg[125]  ( .D(n380), .CLK(clk), .Q(
        decodedPacket1_o[125]) );
  DFFX1 \decodedPacket1_o_reg[124]  ( .D(n379), .CLK(clk), .Q(
        decodedPacket1_o[124]) );
  DFFX1 \decodedPacket1_o_reg[123]  ( .D(n378), .CLK(clk), .Q(
        decodedPacket1_o[123]) );
  DFFX1 \decodedPacket1_o_reg[122]  ( .D(n377), .CLK(clk), .Q(
        decodedPacket1_o[122]) );
  DFFX1 \decodedPacket1_o_reg[121]  ( .D(n376), .CLK(clk), .Q(
        decodedPacket1_o[121]) );
  DFFX1 \decodedPacket1_o_reg[120]  ( .D(n375), .CLK(clk), .Q(
        decodedPacket1_o[120]) );
  DFFX1 \decodedPacket1_o_reg[119]  ( .D(n374), .CLK(clk), .Q(
        decodedPacket1_o[119]) );
  DFFX1 \decodedPacket1_o_reg[118]  ( .D(n373), .CLK(clk), .Q(
        decodedPacket1_o[118]) );
  DFFX1 \decodedPacket1_o_reg[117]  ( .D(n372), .CLK(clk), .Q(
        decodedPacket1_o[117]) );
  DFFX1 \decodedPacket1_o_reg[116]  ( .D(n371), .CLK(clk), .Q(
        decodedPacket1_o[116]) );
  DFFX1 \decodedPacket1_o_reg[115]  ( .D(n370), .CLK(clk), .Q(
        decodedPacket1_o[115]) );
  DFFX1 \decodedPacket1_o_reg[114]  ( .D(n369), .CLK(clk), .Q(
        decodedPacket1_o[114]) );
  DFFX1 \decodedPacket1_o_reg[113]  ( .D(n368), .CLK(clk), .Q(
        decodedPacket1_o[113]) );
  DFFX1 \decodedPacket1_o_reg[112]  ( .D(n367), .CLK(clk), .Q(
        decodedPacket1_o[112]) );
  DFFX1 \decodedPacket1_o_reg[111]  ( .D(n366), .CLK(clk), .Q(
        decodedPacket1_o[111]) );
  DFFX1 \decodedPacket1_o_reg[110]  ( .D(n365), .CLK(clk), .Q(
        decodedPacket1_o[110]) );
  DFFX1 \decodedPacket1_o_reg[109]  ( .D(n364), .CLK(clk), .Q(
        decodedPacket1_o[109]) );
  DFFX1 \decodedPacket1_o_reg[108]  ( .D(n363), .CLK(clk), .Q(
        decodedPacket1_o[108]) );
  DFFX1 \decodedPacket1_o_reg[107]  ( .D(n362), .CLK(clk), .Q(
        decodedPacket1_o[107]) );
  DFFX1 \decodedPacket1_o_reg[106]  ( .D(n361), .CLK(clk), .Q(
        decodedPacket1_o[106]) );
  DFFX1 \decodedPacket1_o_reg[105]  ( .D(n360), .CLK(clk), .Q(
        decodedPacket1_o[105]) );
  DFFX1 \decodedPacket1_o_reg[104]  ( .D(n359), .CLK(clk), .Q(
        decodedPacket1_o[104]) );
  DFFX1 \decodedPacket1_o_reg[103]  ( .D(n358), .CLK(clk), .Q(
        decodedPacket1_o[103]) );
  DFFX1 \decodedPacket1_o_reg[102]  ( .D(n357), .CLK(clk), .Q(
        decodedPacket1_o[102]) );
  DFFX1 \decodedPacket1_o_reg[101]  ( .D(n356), .CLK(clk), .Q(
        decodedPacket1_o[101]) );
  DFFX1 \decodedPacket1_o_reg[100]  ( .D(n355), .CLK(clk), .Q(
        decodedPacket1_o[100]) );
  DFFX1 \decodedPacket1_o_reg[99]  ( .D(n354), .CLK(clk), .Q(
        decodedPacket1_o[99]) );
  DFFX1 \decodedPacket1_o_reg[98]  ( .D(n353), .CLK(clk), .Q(
        decodedPacket1_o[98]) );
  DFFX1 \decodedPacket1_o_reg[97]  ( .D(n352), .CLK(clk), .Q(
        decodedPacket1_o[97]) );
  DFFX1 \decodedPacket1_o_reg[96]  ( .D(n351), .CLK(clk), .Q(
        decodedPacket1_o[96]) );
  DFFX1 \decodedPacket1_o_reg[95]  ( .D(n350), .CLK(clk), .Q(
        decodedPacket1_o[95]) );
  DFFX1 \decodedPacket1_o_reg[94]  ( .D(n349), .CLK(clk), .Q(
        decodedPacket1_o[94]) );
  DFFX1 \decodedPacket1_o_reg[93]  ( .D(n348), .CLK(clk), .Q(
        decodedPacket1_o[93]) );
  DFFX1 \decodedPacket1_o_reg[92]  ( .D(n347), .CLK(clk), .Q(
        decodedPacket1_o[92]) );
  DFFX1 \decodedPacket1_o_reg[91]  ( .D(n346), .CLK(clk), .Q(
        decodedPacket1_o[91]) );
  DFFX1 \decodedPacket1_o_reg[90]  ( .D(n345), .CLK(clk), .Q(
        decodedPacket1_o[90]) );
  DFFX1 \decodedPacket1_o_reg[89]  ( .D(n344), .CLK(clk), .Q(
        decodedPacket1_o[89]) );
  DFFX1 \decodedPacket1_o_reg[88]  ( .D(n343), .CLK(clk), .Q(
        decodedPacket1_o[88]) );
  DFFX1 \decodedPacket1_o_reg[87]  ( .D(n342), .CLK(clk), .Q(
        decodedPacket1_o[87]) );
  DFFX1 \decodedPacket1_o_reg[86]  ( .D(n341), .CLK(clk), .Q(
        decodedPacket1_o[86]) );
  DFFX1 \decodedPacket1_o_reg[85]  ( .D(n340), .CLK(clk), .Q(
        decodedPacket1_o[85]) );
  DFFX1 \decodedPacket1_o_reg[84]  ( .D(n339), .CLK(clk), .Q(
        decodedPacket1_o[84]) );
  DFFX1 \decodedPacket1_o_reg[83]  ( .D(n338), .CLK(clk), .Q(
        decodedPacket1_o[83]) );
  DFFX1 \decodedPacket1_o_reg[82]  ( .D(n337), .CLK(clk), .Q(
        decodedPacket1_o[82]) );
  DFFX1 \decodedPacket1_o_reg[81]  ( .D(n336), .CLK(clk), .Q(
        decodedPacket1_o[81]) );
  DFFX1 \decodedPacket1_o_reg[80]  ( .D(n335), .CLK(clk), .Q(
        decodedPacket1_o[80]) );
  DFFX1 \decodedPacket1_o_reg[79]  ( .D(n334), .CLK(clk), .Q(
        decodedPacket1_o[79]) );
  DFFX1 \decodedPacket1_o_reg[78]  ( .D(n333), .CLK(clk), .Q(
        decodedPacket1_o[78]) );
  DFFX1 \decodedPacket1_o_reg[77]  ( .D(n332), .CLK(clk), .Q(
        decodedPacket1_o[77]) );
  DFFX1 \decodedPacket1_o_reg[76]  ( .D(n331), .CLK(clk), .Q(
        decodedPacket1_o[76]) );
  DFFX1 \decodedPacket1_o_reg[75]  ( .D(n330), .CLK(clk), .Q(
        decodedPacket1_o[75]) );
  DFFX1 \decodedPacket1_o_reg[74]  ( .D(n329), .CLK(clk), .Q(
        decodedPacket1_o[74]) );
  DFFX1 \decodedPacket1_o_reg[73]  ( .D(n328), .CLK(clk), .Q(
        decodedPacket1_o[73]) );
  DFFX1 \decodedPacket1_o_reg[72]  ( .D(n327), .CLK(clk), .Q(
        decodedPacket1_o[72]) );
  DFFX1 \decodedPacket1_o_reg[71]  ( .D(n326), .CLK(clk), .Q(
        decodedPacket1_o[71]) );
  DFFX1 \decodedPacket1_o_reg[70]  ( .D(n325), .CLK(clk), .Q(
        decodedPacket1_o[70]) );
  DFFX1 \decodedPacket1_o_reg[69]  ( .D(n324), .CLK(clk), .Q(
        decodedPacket1_o[69]) );
  DFFX1 \decodedPacket1_o_reg[68]  ( .D(n323), .CLK(clk), .Q(
        decodedPacket1_o[68]) );
  DFFX1 \decodedPacket1_o_reg[67]  ( .D(n322), .CLK(clk), .Q(
        decodedPacket1_o[67]) );
  DFFX1 \decodedPacket1_o_reg[66]  ( .D(n321), .CLK(clk), .Q(
        decodedPacket1_o[66]) );
  DFFX1 \decodedPacket1_o_reg[65]  ( .D(n320), .CLK(clk), .Q(
        decodedPacket1_o[65]) );
  DFFX1 \decodedPacket1_o_reg[64]  ( .D(n319), .CLK(clk), .Q(
        decodedPacket1_o[64]) );
  DFFX1 \decodedPacket1_o_reg[63]  ( .D(n318), .CLK(clk), .Q(
        decodedPacket1_o[63]) );
  DFFX1 \decodedPacket1_o_reg[62]  ( .D(n317), .CLK(clk), .Q(
        decodedPacket1_o[62]) );
  DFFX1 \decodedPacket1_o_reg[61]  ( .D(n316), .CLK(clk), .Q(
        decodedPacket1_o[61]) );
  DFFX1 \decodedPacket1_o_reg[60]  ( .D(n315), .CLK(clk), .Q(
        decodedPacket1_o[60]) );
  DFFX1 \decodedPacket1_o_reg[59]  ( .D(n314), .CLK(clk), .Q(
        decodedPacket1_o[59]) );
  DFFX1 \decodedPacket1_o_reg[58]  ( .D(n313), .CLK(clk), .Q(
        decodedPacket1_o[58]) );
  DFFX1 \decodedPacket1_o_reg[57]  ( .D(n312), .CLK(clk), .Q(
        decodedPacket1_o[57]) );
  DFFX1 \decodedPacket1_o_reg[56]  ( .D(n311), .CLK(clk), .Q(
        decodedPacket1_o[56]) );
  DFFX1 \decodedPacket1_o_reg[55]  ( .D(n310), .CLK(clk), .Q(
        decodedPacket1_o[55]) );
  DFFX1 \decodedPacket1_o_reg[54]  ( .D(n309), .CLK(clk), .Q(
        decodedPacket1_o[54]) );
  DFFX1 \decodedPacket1_o_reg[53]  ( .D(n308), .CLK(clk), .Q(
        decodedPacket1_o[53]) );
  DFFX1 \decodedPacket1_o_reg[52]  ( .D(n307), .CLK(clk), .Q(
        decodedPacket1_o[52]) );
  DFFX1 \decodedPacket1_o_reg[51]  ( .D(n306), .CLK(clk), .Q(
        decodedPacket1_o[51]) );
  DFFX1 \decodedPacket1_o_reg[50]  ( .D(n305), .CLK(clk), .Q(
        decodedPacket1_o[50]) );
  DFFX1 \decodedPacket1_o_reg[49]  ( .D(n304), .CLK(clk), .Q(
        decodedPacket1_o[49]) );
  DFFX1 \decodedPacket1_o_reg[48]  ( .D(n303), .CLK(clk), .Q(
        decodedPacket1_o[48]) );
  DFFX1 \decodedPacket1_o_reg[47]  ( .D(n302), .CLK(clk), .Q(
        decodedPacket1_o[47]) );
  DFFX1 \decodedPacket1_o_reg[46]  ( .D(n301), .CLK(clk), .Q(
        decodedPacket1_o[46]) );
  DFFX1 \decodedPacket1_o_reg[45]  ( .D(n300), .CLK(clk), .Q(
        decodedPacket1_o[45]) );
  DFFX1 \decodedPacket1_o_reg[44]  ( .D(n299), .CLK(clk), .Q(
        decodedPacket1_o[44]) );
  DFFX1 \decodedPacket1_o_reg[43]  ( .D(n298), .CLK(clk), .Q(
        decodedPacket1_o[43]) );
  DFFX1 \decodedPacket1_o_reg[42]  ( .D(n297), .CLK(clk), .Q(
        decodedPacket1_o[42]) );
  DFFX1 \decodedPacket1_o_reg[41]  ( .D(n296), .CLK(clk), .Q(
        decodedPacket1_o[41]) );
  DFFX1 \decodedPacket1_o_reg[40]  ( .D(n295), .CLK(clk), .Q(
        decodedPacket1_o[40]) );
  DFFX1 \decodedPacket1_o_reg[39]  ( .D(n294), .CLK(clk), .Q(
        decodedPacket1_o[39]) );
  DFFX1 \decodedPacket1_o_reg[38]  ( .D(n293), .CLK(clk), .Q(
        decodedPacket1_o[38]) );
  DFFX1 \decodedPacket1_o_reg[37]  ( .D(n292), .CLK(clk), .Q(
        decodedPacket1_o[37]) );
  DFFX1 \decodedPacket1_o_reg[36]  ( .D(n291), .CLK(clk), .Q(
        decodedPacket1_o[36]) );
  DFFX1 \decodedPacket1_o_reg[35]  ( .D(n290), .CLK(clk), .Q(
        decodedPacket1_o[35]) );
  DFFX1 \decodedPacket1_o_reg[34]  ( .D(n289), .CLK(clk), .Q(
        decodedPacket1_o[34]) );
  DFFX1 \decodedPacket1_o_reg[33]  ( .D(n288), .CLK(clk), .Q(
        decodedPacket1_o[33]) );
  DFFX1 \decodedPacket1_o_reg[32]  ( .D(n287), .CLK(clk), .Q(
        decodedPacket1_o[32]) );
  DFFX1 \decodedPacket1_o_reg[31]  ( .D(n286), .CLK(clk), .Q(
        decodedPacket1_o[31]) );
  DFFX1 \decodedPacket1_o_reg[30]  ( .D(n285), .CLK(clk), .Q(
        decodedPacket1_o[30]) );
  DFFX1 \decodedPacket1_o_reg[29]  ( .D(n284), .CLK(clk), .Q(
        decodedPacket1_o[29]) );
  DFFX1 \decodedPacket1_o_reg[28]  ( .D(n283), .CLK(clk), .Q(
        decodedPacket1_o[28]) );
  DFFX1 \decodedPacket1_o_reg[27]  ( .D(n282), .CLK(clk), .Q(
        decodedPacket1_o[27]) );
  DFFX1 \decodedPacket1_o_reg[26]  ( .D(n281), .CLK(clk), .Q(
        decodedPacket1_o[26]) );
  DFFX1 \decodedPacket1_o_reg[25]  ( .D(n280), .CLK(clk), .Q(
        decodedPacket1_o[25]) );
  DFFX1 \decodedPacket1_o_reg[24]  ( .D(n279), .CLK(clk), .Q(
        decodedPacket1_o[24]) );
  DFFX1 \decodedPacket1_o_reg[23]  ( .D(n278), .CLK(clk), .Q(
        decodedPacket1_o[23]) );
  DFFX1 \decodedPacket1_o_reg[22]  ( .D(n277), .CLK(clk), .Q(
        decodedPacket1_o[22]) );
  DFFX1 \decodedPacket1_o_reg[21]  ( .D(n276), .CLK(clk), .Q(
        decodedPacket1_o[21]) );
  DFFX1 \decodedPacket1_o_reg[20]  ( .D(n275), .CLK(clk), .Q(
        decodedPacket1_o[20]) );
  DFFX1 \decodedPacket1_o_reg[19]  ( .D(n274), .CLK(clk), .Q(
        decodedPacket1_o[19]) );
  DFFX1 \decodedPacket1_o_reg[18]  ( .D(n273), .CLK(clk), .Q(
        decodedPacket1_o[18]) );
  DFFX1 \decodedPacket1_o_reg[17]  ( .D(n272), .CLK(clk), .Q(
        decodedPacket1_o[17]) );
  DFFX1 \decodedPacket1_o_reg[16]  ( .D(n271), .CLK(clk), .Q(
        decodedPacket1_o[16]) );
  DFFX1 \decodedPacket1_o_reg[15]  ( .D(n270), .CLK(clk), .Q(
        decodedPacket1_o[15]) );
  DFFX1 \decodedPacket1_o_reg[14]  ( .D(n269), .CLK(clk), .Q(
        decodedPacket1_o[14]) );
  DFFX1 \decodedPacket1_o_reg[13]  ( .D(n268), .CLK(clk), .Q(
        decodedPacket1_o[13]) );
  DFFX1 \decodedPacket1_o_reg[12]  ( .D(n267), .CLK(clk), .Q(
        decodedPacket1_o[12]) );
  DFFX1 \decodedPacket1_o_reg[11]  ( .D(n266), .CLK(clk), .Q(
        decodedPacket1_o[11]) );
  DFFX1 \decodedPacket1_o_reg[10]  ( .D(n265), .CLK(clk), .Q(
        decodedPacket1_o[10]) );
  DFFX1 \decodedPacket1_o_reg[9]  ( .D(n264), .CLK(clk), .Q(
        decodedPacket1_o[9]) );
  DFFX1 \decodedPacket1_o_reg[8]  ( .D(n263), .CLK(clk), .Q(
        decodedPacket1_o[8]) );
  DFFX1 \decodedPacket1_o_reg[7]  ( .D(n262), .CLK(clk), .Q(
        decodedPacket1_o[7]) );
  DFFX1 \decodedPacket1_o_reg[6]  ( .D(n261), .CLK(clk), .Q(
        decodedPacket1_o[6]) );
  DFFX1 \decodedPacket1_o_reg[5]  ( .D(n260), .CLK(clk), .Q(
        decodedPacket1_o[5]) );
  DFFX1 \decodedPacket1_o_reg[4]  ( .D(n259), .CLK(clk), .Q(
        decodedPacket1_o[4]) );
  DFFX1 \decodedPacket1_o_reg[3]  ( .D(n258), .CLK(clk), .Q(
        decodedPacket1_o[3]) );
  DFFX1 \decodedPacket1_o_reg[2]  ( .D(n257), .CLK(clk), .Q(
        decodedPacket1_o[2]) );
  DFFX1 \decodedPacket1_o_reg[1]  ( .D(n256), .CLK(clk), .Q(
        decodedPacket1_o[1]) );
  DFFX1 \decodedPacket1_o_reg[0]  ( .D(n255), .CLK(clk), .Q(
        decodedPacket1_o[0]) );
  DFFX1 \decodedPacket2_o_reg[125]  ( .D(n254), .CLK(clk), .Q(
        decodedPacket2_o[125]) );
  DFFX1 \decodedPacket2_o_reg[124]  ( .D(n253), .CLK(clk), .Q(
        decodedPacket2_o[124]) );
  DFFX1 \decodedPacket2_o_reg[123]  ( .D(n252), .CLK(clk), .Q(
        decodedPacket2_o[123]) );
  DFFX1 \decodedPacket2_o_reg[122]  ( .D(n251), .CLK(clk), .Q(
        decodedPacket2_o[122]) );
  DFFX1 \decodedPacket2_o_reg[121]  ( .D(n250), .CLK(clk), .Q(
        decodedPacket2_o[121]) );
  DFFX1 \decodedPacket2_o_reg[120]  ( .D(n249), .CLK(clk), .Q(
        decodedPacket2_o[120]) );
  DFFX1 \decodedPacket2_o_reg[119]  ( .D(n248), .CLK(clk), .Q(
        decodedPacket2_o[119]) );
  DFFX1 \decodedPacket2_o_reg[118]  ( .D(n247), .CLK(clk), .Q(
        decodedPacket2_o[118]) );
  DFFX1 \decodedPacket2_o_reg[117]  ( .D(n246), .CLK(clk), .Q(
        decodedPacket2_o[117]) );
  DFFX1 \decodedPacket2_o_reg[116]  ( .D(n245), .CLK(clk), .Q(
        decodedPacket2_o[116]) );
  DFFX1 \decodedPacket2_o_reg[115]  ( .D(n244), .CLK(clk), .Q(
        decodedPacket2_o[115]) );
  DFFX1 \decodedPacket2_o_reg[114]  ( .D(n243), .CLK(clk), .Q(
        decodedPacket2_o[114]) );
  DFFX1 \decodedPacket2_o_reg[113]  ( .D(n242), .CLK(clk), .Q(
        decodedPacket2_o[113]) );
  DFFX1 \decodedPacket2_o_reg[112]  ( .D(n241), .CLK(clk), .Q(
        decodedPacket2_o[112]) );
  DFFX1 \decodedPacket2_o_reg[111]  ( .D(n240), .CLK(clk), .Q(
        decodedPacket2_o[111]) );
  DFFX1 \decodedPacket2_o_reg[110]  ( .D(n239), .CLK(clk), .Q(
        decodedPacket2_o[110]) );
  DFFX1 \decodedPacket2_o_reg[109]  ( .D(n238), .CLK(clk), .Q(
        decodedPacket2_o[109]) );
  DFFX1 \decodedPacket2_o_reg[108]  ( .D(n237), .CLK(clk), .Q(
        decodedPacket2_o[108]) );
  DFFX1 \decodedPacket2_o_reg[107]  ( .D(n236), .CLK(clk), .Q(
        decodedPacket2_o[107]) );
  DFFX1 \decodedPacket2_o_reg[106]  ( .D(n235), .CLK(clk), .Q(
        decodedPacket2_o[106]) );
  DFFX1 \decodedPacket2_o_reg[105]  ( .D(n234), .CLK(clk), .Q(
        decodedPacket2_o[105]) );
  DFFX1 \decodedPacket2_o_reg[104]  ( .D(n233), .CLK(clk), .Q(
        decodedPacket2_o[104]) );
  DFFX1 \decodedPacket2_o_reg[103]  ( .D(n232), .CLK(clk), .Q(
        decodedPacket2_o[103]) );
  DFFX1 \decodedPacket2_o_reg[102]  ( .D(n231), .CLK(clk), .Q(
        decodedPacket2_o[102]) );
  DFFX1 \decodedPacket2_o_reg[101]  ( .D(n230), .CLK(clk), .Q(
        decodedPacket2_o[101]) );
  DFFX1 \decodedPacket2_o_reg[100]  ( .D(n229), .CLK(clk), .Q(
        decodedPacket2_o[100]) );
  DFFX1 \decodedPacket2_o_reg[99]  ( .D(n228), .CLK(clk), .Q(
        decodedPacket2_o[99]) );
  DFFX1 \decodedPacket2_o_reg[98]  ( .D(n227), .CLK(clk), .Q(
        decodedPacket2_o[98]) );
  DFFX1 \decodedPacket2_o_reg[97]  ( .D(n226), .CLK(clk), .Q(
        decodedPacket2_o[97]) );
  DFFX1 \decodedPacket2_o_reg[96]  ( .D(n225), .CLK(clk), .Q(
        decodedPacket2_o[96]) );
  DFFX1 \decodedPacket2_o_reg[95]  ( .D(n224), .CLK(clk), .Q(
        decodedPacket2_o[95]) );
  DFFX1 \decodedPacket2_o_reg[94]  ( .D(n223), .CLK(clk), .Q(
        decodedPacket2_o[94]) );
  DFFX1 \decodedPacket2_o_reg[93]  ( .D(n222), .CLK(clk), .Q(
        decodedPacket2_o[93]) );
  DFFX1 \decodedPacket2_o_reg[92]  ( .D(n221), .CLK(clk), .Q(
        decodedPacket2_o[92]) );
  DFFX1 \decodedPacket2_o_reg[91]  ( .D(n220), .CLK(clk), .Q(
        decodedPacket2_o[91]) );
  DFFX1 \decodedPacket2_o_reg[90]  ( .D(n219), .CLK(clk), .Q(
        decodedPacket2_o[90]) );
  DFFX1 \decodedPacket2_o_reg[89]  ( .D(n218), .CLK(clk), .Q(
        decodedPacket2_o[89]) );
  DFFX1 \decodedPacket2_o_reg[88]  ( .D(n217), .CLK(clk), .Q(
        decodedPacket2_o[88]) );
  DFFX1 \decodedPacket2_o_reg[87]  ( .D(n216), .CLK(clk), .Q(
        decodedPacket2_o[87]) );
  DFFX1 \decodedPacket2_o_reg[86]  ( .D(n215), .CLK(clk), .Q(
        decodedPacket2_o[86]) );
  DFFX1 \decodedPacket2_o_reg[85]  ( .D(n214), .CLK(clk), .Q(
        decodedPacket2_o[85]) );
  DFFX1 \decodedPacket2_o_reg[84]  ( .D(n213), .CLK(clk), .Q(
        decodedPacket2_o[84]) );
  DFFX1 \decodedPacket2_o_reg[83]  ( .D(n212), .CLK(clk), .Q(
        decodedPacket2_o[83]) );
  DFFX1 \decodedPacket2_o_reg[82]  ( .D(n211), .CLK(clk), .Q(
        decodedPacket2_o[82]) );
  DFFX1 \decodedPacket2_o_reg[81]  ( .D(n210), .CLK(clk), .Q(
        decodedPacket2_o[81]) );
  DFFX1 \decodedPacket2_o_reg[80]  ( .D(n209), .CLK(clk), .Q(
        decodedPacket2_o[80]) );
  DFFX1 \decodedPacket2_o_reg[79]  ( .D(n208), .CLK(clk), .Q(
        decodedPacket2_o[79]) );
  DFFX1 \decodedPacket2_o_reg[78]  ( .D(n207), .CLK(clk), .Q(
        decodedPacket2_o[78]) );
  DFFX1 \decodedPacket2_o_reg[77]  ( .D(n206), .CLK(clk), .Q(
        decodedPacket2_o[77]) );
  DFFX1 \decodedPacket2_o_reg[76]  ( .D(n205), .CLK(clk), .Q(
        decodedPacket2_o[76]) );
  DFFX1 \decodedPacket2_o_reg[75]  ( .D(n204), .CLK(clk), .Q(
        decodedPacket2_o[75]) );
  DFFX1 \decodedPacket2_o_reg[74]  ( .D(n203), .CLK(clk), .Q(
        decodedPacket2_o[74]) );
  DFFX1 \decodedPacket2_o_reg[73]  ( .D(n202), .CLK(clk), .Q(
        decodedPacket2_o[73]) );
  DFFX1 \decodedPacket2_o_reg[72]  ( .D(n201), .CLK(clk), .Q(
        decodedPacket2_o[72]) );
  DFFX1 \decodedPacket2_o_reg[71]  ( .D(n200), .CLK(clk), .Q(
        decodedPacket2_o[71]) );
  DFFX1 \decodedPacket2_o_reg[70]  ( .D(n199), .CLK(clk), .Q(
        decodedPacket2_o[70]) );
  DFFX1 \decodedPacket2_o_reg[69]  ( .D(n198), .CLK(clk), .Q(
        decodedPacket2_o[69]) );
  DFFX1 \decodedPacket2_o_reg[68]  ( .D(n197), .CLK(clk), .Q(
        decodedPacket2_o[68]) );
  DFFX1 \decodedPacket2_o_reg[67]  ( .D(n196), .CLK(clk), .Q(
        decodedPacket2_o[67]) );
  DFFX1 \decodedPacket2_o_reg[66]  ( .D(n195), .CLK(clk), .Q(
        decodedPacket2_o[66]) );
  DFFX1 \decodedPacket2_o_reg[65]  ( .D(n194), .CLK(clk), .Q(
        decodedPacket2_o[65]) );
  DFFX1 \decodedPacket2_o_reg[64]  ( .D(n193), .CLK(clk), .Q(
        decodedPacket2_o[64]) );
  DFFX1 \decodedPacket2_o_reg[63]  ( .D(n192), .CLK(clk), .Q(
        decodedPacket2_o[63]) );
  DFFX1 \decodedPacket2_o_reg[62]  ( .D(n191), .CLK(clk), .Q(
        decodedPacket2_o[62]) );
  DFFX1 \decodedPacket2_o_reg[61]  ( .D(n190), .CLK(clk), .Q(
        decodedPacket2_o[61]) );
  DFFX1 \decodedPacket2_o_reg[60]  ( .D(n189), .CLK(clk), .Q(
        decodedPacket2_o[60]) );
  DFFX1 \decodedPacket2_o_reg[59]  ( .D(n188), .CLK(clk), .Q(
        decodedPacket2_o[59]) );
  DFFX1 \decodedPacket2_o_reg[58]  ( .D(n187), .CLK(clk), .Q(
        decodedPacket2_o[58]) );
  DFFX1 \decodedPacket2_o_reg[57]  ( .D(n186), .CLK(clk), .Q(
        decodedPacket2_o[57]) );
  DFFX1 \decodedPacket2_o_reg[56]  ( .D(n185), .CLK(clk), .Q(
        decodedPacket2_o[56]) );
  DFFX1 \decodedPacket2_o_reg[55]  ( .D(n184), .CLK(clk), .Q(
        decodedPacket2_o[55]) );
  DFFX1 \decodedPacket2_o_reg[54]  ( .D(n183), .CLK(clk), .Q(
        decodedPacket2_o[54]) );
  DFFX1 \decodedPacket2_o_reg[53]  ( .D(n182), .CLK(clk), .Q(
        decodedPacket2_o[53]) );
  DFFX1 \decodedPacket2_o_reg[52]  ( .D(n181), .CLK(clk), .Q(
        decodedPacket2_o[52]) );
  DFFX1 \decodedPacket2_o_reg[51]  ( .D(n180), .CLK(clk), .Q(
        decodedPacket2_o[51]) );
  DFFX1 \decodedPacket2_o_reg[50]  ( .D(n179), .CLK(clk), .Q(
        decodedPacket2_o[50]) );
  DFFX1 \decodedPacket2_o_reg[49]  ( .D(n178), .CLK(clk), .Q(
        decodedPacket2_o[49]) );
  DFFX1 \decodedPacket2_o_reg[48]  ( .D(n177), .CLK(clk), .Q(
        decodedPacket2_o[48]) );
  DFFX1 \decodedPacket2_o_reg[47]  ( .D(n176), .CLK(clk), .Q(
        decodedPacket2_o[47]) );
  DFFX1 \decodedPacket2_o_reg[46]  ( .D(n175), .CLK(clk), .Q(
        decodedPacket2_o[46]) );
  DFFX1 \decodedPacket2_o_reg[45]  ( .D(n174), .CLK(clk), .Q(
        decodedPacket2_o[45]) );
  DFFX1 \decodedPacket2_o_reg[44]  ( .D(n173), .CLK(clk), .Q(
        decodedPacket2_o[44]) );
  DFFX1 \decodedPacket2_o_reg[43]  ( .D(n172), .CLK(clk), .Q(
        decodedPacket2_o[43]) );
  DFFX1 \decodedPacket2_o_reg[42]  ( .D(n171), .CLK(clk), .Q(
        decodedPacket2_o[42]) );
  DFFX1 \decodedPacket2_o_reg[41]  ( .D(n170), .CLK(clk), .Q(
        decodedPacket2_o[41]) );
  DFFX1 \decodedPacket2_o_reg[40]  ( .D(n169), .CLK(clk), .Q(
        decodedPacket2_o[40]) );
  DFFX1 \decodedPacket2_o_reg[39]  ( .D(n168), .CLK(clk), .Q(
        decodedPacket2_o[39]) );
  DFFX1 \decodedPacket2_o_reg[38]  ( .D(n167), .CLK(clk), .Q(
        decodedPacket2_o[38]) );
  DFFX1 \decodedPacket2_o_reg[37]  ( .D(n166), .CLK(clk), .Q(
        decodedPacket2_o[37]) );
  DFFX1 \decodedPacket2_o_reg[36]  ( .D(n165), .CLK(clk), .Q(
        decodedPacket2_o[36]) );
  DFFX1 \decodedPacket2_o_reg[35]  ( .D(n164), .CLK(clk), .Q(
        decodedPacket2_o[35]) );
  DFFX1 \decodedPacket2_o_reg[34]  ( .D(n163), .CLK(clk), .Q(
        decodedPacket2_o[34]) );
  DFFX1 \decodedPacket2_o_reg[33]  ( .D(n162), .CLK(clk), .Q(
        decodedPacket2_o[33]) );
  DFFX1 \decodedPacket2_o_reg[32]  ( .D(n161), .CLK(clk), .Q(
        decodedPacket2_o[32]) );
  DFFX1 \decodedPacket2_o_reg[31]  ( .D(n160), .CLK(clk), .Q(
        decodedPacket2_o[31]) );
  DFFX1 \decodedPacket2_o_reg[30]  ( .D(n159), .CLK(clk), .Q(
        decodedPacket2_o[30]) );
  DFFX1 \decodedPacket2_o_reg[29]  ( .D(n158), .CLK(clk), .Q(
        decodedPacket2_o[29]) );
  DFFX1 \decodedPacket2_o_reg[28]  ( .D(n157), .CLK(clk), .Q(
        decodedPacket2_o[28]) );
  DFFX1 \decodedPacket2_o_reg[27]  ( .D(n156), .CLK(clk), .Q(
        decodedPacket2_o[27]) );
  DFFX1 \decodedPacket2_o_reg[26]  ( .D(n155), .CLK(clk), .Q(
        decodedPacket2_o[26]) );
  DFFX1 \decodedPacket2_o_reg[25]  ( .D(n154), .CLK(clk), .Q(
        decodedPacket2_o[25]) );
  DFFX1 \decodedPacket2_o_reg[24]  ( .D(n153), .CLK(clk), .Q(
        decodedPacket2_o[24]) );
  DFFX1 \decodedPacket2_o_reg[23]  ( .D(n152), .CLK(clk), .Q(
        decodedPacket2_o[23]) );
  DFFX1 \decodedPacket2_o_reg[22]  ( .D(n151), .CLK(clk), .Q(
        decodedPacket2_o[22]) );
  DFFX1 \decodedPacket2_o_reg[21]  ( .D(n150), .CLK(clk), .Q(
        decodedPacket2_o[21]) );
  DFFX1 \decodedPacket2_o_reg[20]  ( .D(n149), .CLK(clk), .Q(
        decodedPacket2_o[20]) );
  DFFX1 \decodedPacket2_o_reg[19]  ( .D(n148), .CLK(clk), .Q(
        decodedPacket2_o[19]) );
  DFFX1 \decodedPacket2_o_reg[18]  ( .D(n147), .CLK(clk), .Q(
        decodedPacket2_o[18]) );
  DFFX1 \decodedPacket2_o_reg[17]  ( .D(n146), .CLK(clk), .Q(
        decodedPacket2_o[17]) );
  DFFX1 \decodedPacket2_o_reg[16]  ( .D(n145), .CLK(clk), .Q(
        decodedPacket2_o[16]) );
  DFFX1 \decodedPacket2_o_reg[15]  ( .D(n144), .CLK(clk), .Q(
        decodedPacket2_o[15]) );
  DFFX1 \decodedPacket2_o_reg[14]  ( .D(n143), .CLK(clk), .Q(
        decodedPacket2_o[14]) );
  DFFX1 \decodedPacket2_o_reg[13]  ( .D(n142), .CLK(clk), .Q(
        decodedPacket2_o[13]) );
  DFFX1 \decodedPacket2_o_reg[12]  ( .D(n141), .CLK(clk), .Q(
        decodedPacket2_o[12]) );
  DFFX1 \decodedPacket2_o_reg[11]  ( .D(n140), .CLK(clk), .Q(
        decodedPacket2_o[11]) );
  DFFX1 \decodedPacket2_o_reg[10]  ( .D(n139), .CLK(clk), .Q(
        decodedPacket2_o[10]) );
  DFFX1 \decodedPacket2_o_reg[9]  ( .D(n138), .CLK(clk), .Q(
        decodedPacket2_o[9]) );
  DFFX1 \decodedPacket2_o_reg[8]  ( .D(n137), .CLK(clk), .Q(
        decodedPacket2_o[8]) );
  DFFX1 \decodedPacket2_o_reg[7]  ( .D(n136), .CLK(clk), .Q(
        decodedPacket2_o[7]) );
  DFFX1 \decodedPacket2_o_reg[6]  ( .D(n135), .CLK(clk), .Q(
        decodedPacket2_o[6]) );
  DFFX1 \decodedPacket2_o_reg[5]  ( .D(n134), .CLK(clk), .Q(
        decodedPacket2_o[5]) );
  DFFX1 \decodedPacket2_o_reg[4]  ( .D(n133), .CLK(clk), .Q(
        decodedPacket2_o[4]) );
  DFFX1 \decodedPacket2_o_reg[3]  ( .D(n132), .CLK(clk), .Q(
        decodedPacket2_o[3]) );
  DFFX1 \decodedPacket2_o_reg[2]  ( .D(n131), .CLK(clk), .Q(
        decodedPacket2_o[2]) );
  DFFX1 \decodedPacket2_o_reg[1]  ( .D(n130), .CLK(clk), .Q(
        decodedPacket2_o[1]) );
  DFFX1 \decodedPacket2_o_reg[0]  ( .D(n129), .CLK(clk), .Q(
        decodedPacket2_o[0]) );
  DFFX1 \decodedPacket3_o_reg[125]  ( .D(n128), .CLK(clk), .Q(
        decodedPacket3_o[125]) );
  DFFX1 \decodedPacket3_o_reg[124]  ( .D(n127), .CLK(clk), .Q(
        decodedPacket3_o[124]) );
  DFFX1 \decodedPacket3_o_reg[123]  ( .D(n126), .CLK(clk), .Q(
        decodedPacket3_o[123]) );
  DFFX1 \decodedPacket3_o_reg[122]  ( .D(n125), .CLK(clk), .Q(
        decodedPacket3_o[122]) );
  DFFX1 \decodedPacket3_o_reg[121]  ( .D(n124), .CLK(clk), .Q(
        decodedPacket3_o[121]) );
  DFFX1 \decodedPacket3_o_reg[120]  ( .D(n123), .CLK(clk), .Q(
        decodedPacket3_o[120]) );
  DFFX1 \decodedPacket3_o_reg[119]  ( .D(n122), .CLK(clk), .Q(
        decodedPacket3_o[119]) );
  DFFX1 \decodedPacket3_o_reg[118]  ( .D(n121), .CLK(clk), .Q(
        decodedPacket3_o[118]) );
  DFFX1 \decodedPacket3_o_reg[117]  ( .D(n120), .CLK(clk), .Q(
        decodedPacket3_o[117]) );
  DFFX1 \decodedPacket3_o_reg[116]  ( .D(n119), .CLK(clk), .Q(
        decodedPacket3_o[116]) );
  DFFX1 \decodedPacket3_o_reg[115]  ( .D(n118), .CLK(clk), .Q(
        decodedPacket3_o[115]) );
  DFFX1 \decodedPacket3_o_reg[114]  ( .D(n117), .CLK(clk), .Q(
        decodedPacket3_o[114]) );
  DFFX1 \decodedPacket3_o_reg[113]  ( .D(n116), .CLK(clk), .Q(
        decodedPacket3_o[113]) );
  DFFX1 \decodedPacket3_o_reg[112]  ( .D(n115), .CLK(clk), .Q(
        decodedPacket3_o[112]) );
  DFFX1 \decodedPacket3_o_reg[111]  ( .D(n114), .CLK(clk), .Q(
        decodedPacket3_o[111]) );
  DFFX1 \decodedPacket3_o_reg[110]  ( .D(n113), .CLK(clk), .Q(
        decodedPacket3_o[110]) );
  DFFX1 \decodedPacket3_o_reg[109]  ( .D(n112), .CLK(clk), .Q(
        decodedPacket3_o[109]) );
  DFFX1 \decodedPacket3_o_reg[108]  ( .D(n111), .CLK(clk), .Q(
        decodedPacket3_o[108]) );
  DFFX1 \decodedPacket3_o_reg[107]  ( .D(n110), .CLK(clk), .Q(
        decodedPacket3_o[107]) );
  DFFX1 \decodedPacket3_o_reg[106]  ( .D(n109), .CLK(clk), .Q(
        decodedPacket3_o[106]) );
  DFFX1 \decodedPacket3_o_reg[105]  ( .D(n108), .CLK(clk), .Q(
        decodedPacket3_o[105]) );
  DFFX1 \decodedPacket3_o_reg[104]  ( .D(n107), .CLK(clk), .Q(
        decodedPacket3_o[104]) );
  DFFX1 \decodedPacket3_o_reg[103]  ( .D(n106), .CLK(clk), .Q(
        decodedPacket3_o[103]) );
  DFFX1 \decodedPacket3_o_reg[102]  ( .D(n105), .CLK(clk), .Q(
        decodedPacket3_o[102]) );
  DFFX1 \decodedPacket3_o_reg[101]  ( .D(n104), .CLK(clk), .Q(
        decodedPacket3_o[101]) );
  DFFX1 \decodedPacket3_o_reg[100]  ( .D(n103), .CLK(clk), .Q(
        decodedPacket3_o[100]) );
  DFFX1 \decodedPacket3_o_reg[99]  ( .D(n102), .CLK(clk), .Q(
        decodedPacket3_o[99]) );
  DFFX1 \decodedPacket3_o_reg[98]  ( .D(n101), .CLK(clk), .Q(
        decodedPacket3_o[98]) );
  DFFX1 \decodedPacket3_o_reg[97]  ( .D(n100), .CLK(clk), .Q(
        decodedPacket3_o[97]) );
  DFFX1 \decodedPacket3_o_reg[96]  ( .D(n99), .CLK(clk), .Q(
        decodedPacket3_o[96]) );
  DFFX1 \decodedPacket3_o_reg[95]  ( .D(n98), .CLK(clk), .Q(
        decodedPacket3_o[95]) );
  DFFX1 \decodedPacket3_o_reg[94]  ( .D(n97), .CLK(clk), .Q(
        decodedPacket3_o[94]) );
  DFFX1 \decodedPacket3_o_reg[93]  ( .D(n96), .CLK(clk), .Q(
        decodedPacket3_o[93]) );
  DFFX1 \decodedPacket3_o_reg[92]  ( .D(n95), .CLK(clk), .Q(
        decodedPacket3_o[92]) );
  DFFX1 \decodedPacket3_o_reg[91]  ( .D(n94), .CLK(clk), .Q(
        decodedPacket3_o[91]) );
  DFFX1 \decodedPacket3_o_reg[90]  ( .D(n93), .CLK(clk), .Q(
        decodedPacket3_o[90]) );
  DFFX1 \decodedPacket3_o_reg[89]  ( .D(n92), .CLK(clk), .Q(
        decodedPacket3_o[89]) );
  DFFX1 \decodedPacket3_o_reg[88]  ( .D(n91), .CLK(clk), .Q(
        decodedPacket3_o[88]) );
  DFFX1 \decodedPacket3_o_reg[87]  ( .D(n90), .CLK(clk), .Q(
        decodedPacket3_o[87]) );
  DFFX1 \decodedPacket3_o_reg[86]  ( .D(n89), .CLK(clk), .Q(
        decodedPacket3_o[86]) );
  DFFX1 \decodedPacket3_o_reg[85]  ( .D(n88), .CLK(clk), .Q(
        decodedPacket3_o[85]) );
  DFFX1 \decodedPacket3_o_reg[84]  ( .D(n87), .CLK(clk), .Q(
        decodedPacket3_o[84]) );
  DFFX1 \decodedPacket3_o_reg[83]  ( .D(n86), .CLK(clk), .Q(
        decodedPacket3_o[83]) );
  DFFX1 \decodedPacket3_o_reg[82]  ( .D(n85), .CLK(clk), .Q(
        decodedPacket3_o[82]) );
  DFFX1 \decodedPacket3_o_reg[81]  ( .D(n84), .CLK(clk), .Q(
        decodedPacket3_o[81]) );
  DFFX1 \decodedPacket3_o_reg[80]  ( .D(n83), .CLK(clk), .Q(
        decodedPacket3_o[80]) );
  DFFX1 \decodedPacket3_o_reg[79]  ( .D(n82), .CLK(clk), .Q(
        decodedPacket3_o[79]) );
  DFFX1 \decodedPacket3_o_reg[78]  ( .D(n81), .CLK(clk), .Q(
        decodedPacket3_o[78]) );
  DFFX1 \decodedPacket3_o_reg[77]  ( .D(n80), .CLK(clk), .Q(
        decodedPacket3_o[77]) );
  DFFX1 \decodedPacket3_o_reg[76]  ( .D(n79), .CLK(clk), .Q(
        decodedPacket3_o[76]) );
  DFFX1 \decodedPacket3_o_reg[75]  ( .D(n78), .CLK(clk), .Q(
        decodedPacket3_o[75]) );
  DFFX1 \decodedPacket3_o_reg[74]  ( .D(n77), .CLK(clk), .Q(
        decodedPacket3_o[74]) );
  DFFX1 \decodedPacket3_o_reg[73]  ( .D(n76), .CLK(clk), .Q(
        decodedPacket3_o[73]) );
  DFFX1 \decodedPacket3_o_reg[72]  ( .D(n75), .CLK(clk), .Q(
        decodedPacket3_o[72]) );
  DFFX1 \decodedPacket3_o_reg[71]  ( .D(n74), .CLK(clk), .Q(
        decodedPacket3_o[71]) );
  DFFX1 \decodedPacket3_o_reg[70]  ( .D(n73), .CLK(clk), .Q(
        decodedPacket3_o[70]) );
  DFFX1 \decodedPacket3_o_reg[69]  ( .D(n72), .CLK(clk), .Q(
        decodedPacket3_o[69]) );
  DFFX1 \decodedPacket3_o_reg[68]  ( .D(n71), .CLK(clk), .Q(
        decodedPacket3_o[68]) );
  DFFX1 \decodedPacket3_o_reg[67]  ( .D(n70), .CLK(clk), .Q(
        decodedPacket3_o[67]) );
  DFFX1 \decodedPacket3_o_reg[66]  ( .D(n69), .CLK(clk), .Q(
        decodedPacket3_o[66]) );
  DFFX1 \decodedPacket3_o_reg[65]  ( .D(n68), .CLK(clk), .Q(
        decodedPacket3_o[65]) );
  DFFX1 \decodedPacket3_o_reg[64]  ( .D(n67), .CLK(clk), .Q(
        decodedPacket3_o[64]) );
  DFFX1 \decodedPacket3_o_reg[63]  ( .D(n66), .CLK(clk), .Q(
        decodedPacket3_o[63]) );
  DFFX1 \decodedPacket3_o_reg[62]  ( .D(n65), .CLK(clk), .Q(
        decodedPacket3_o[62]) );
  DFFX1 \decodedPacket3_o_reg[61]  ( .D(n64), .CLK(clk), .Q(
        decodedPacket3_o[61]) );
  DFFX1 \decodedPacket3_o_reg[60]  ( .D(n63), .CLK(clk), .Q(
        decodedPacket3_o[60]) );
  DFFX1 \decodedPacket3_o_reg[59]  ( .D(n62), .CLK(clk), .Q(
        decodedPacket3_o[59]) );
  DFFX1 \decodedPacket3_o_reg[58]  ( .D(n61), .CLK(clk), .Q(
        decodedPacket3_o[58]) );
  DFFX1 \decodedPacket3_o_reg[57]  ( .D(n60), .CLK(clk), .Q(
        decodedPacket3_o[57]) );
  DFFX1 \decodedPacket3_o_reg[56]  ( .D(n59), .CLK(clk), .Q(
        decodedPacket3_o[56]) );
  DFFX1 \decodedPacket3_o_reg[55]  ( .D(n58), .CLK(clk), .Q(
        decodedPacket3_o[55]) );
  DFFX1 \decodedPacket3_o_reg[54]  ( .D(n57), .CLK(clk), .Q(
        decodedPacket3_o[54]) );
  DFFX1 \decodedPacket3_o_reg[53]  ( .D(n56), .CLK(clk), .Q(
        decodedPacket3_o[53]) );
  DFFX1 \decodedPacket3_o_reg[52]  ( .D(n55), .CLK(clk), .Q(
        decodedPacket3_o[52]) );
  DFFX1 \decodedPacket3_o_reg[51]  ( .D(n54), .CLK(clk), .Q(
        decodedPacket3_o[51]) );
  DFFX1 \decodedPacket3_o_reg[50]  ( .D(n53), .CLK(clk), .Q(
        decodedPacket3_o[50]) );
  DFFX1 \decodedPacket3_o_reg[49]  ( .D(n52), .CLK(clk), .Q(
        decodedPacket3_o[49]) );
  DFFX1 \decodedPacket3_o_reg[48]  ( .D(n51), .CLK(clk), .Q(
        decodedPacket3_o[48]) );
  DFFX1 \decodedPacket3_o_reg[47]  ( .D(n50), .CLK(clk), .Q(
        decodedPacket3_o[47]) );
  DFFX1 \decodedPacket3_o_reg[46]  ( .D(n49), .CLK(clk), .Q(
        decodedPacket3_o[46]) );
  DFFX1 \decodedPacket3_o_reg[45]  ( .D(n48), .CLK(clk), .Q(
        decodedPacket3_o[45]) );
  DFFX1 \decodedPacket3_o_reg[44]  ( .D(n47), .CLK(clk), .Q(
        decodedPacket3_o[44]) );
  DFFX1 \decodedPacket3_o_reg[43]  ( .D(n46), .CLK(clk), .Q(
        decodedPacket3_o[43]) );
  DFFX1 \decodedPacket3_o_reg[42]  ( .D(n45), .CLK(clk), .Q(
        decodedPacket3_o[42]) );
  DFFX1 \decodedPacket3_o_reg[41]  ( .D(n44), .CLK(clk), .Q(
        decodedPacket3_o[41]) );
  DFFX1 \decodedPacket3_o_reg[40]  ( .D(n43), .CLK(clk), .Q(
        decodedPacket3_o[40]) );
  DFFX1 \decodedPacket3_o_reg[39]  ( .D(n42), .CLK(clk), .Q(
        decodedPacket3_o[39]) );
  DFFX1 \decodedPacket3_o_reg[38]  ( .D(n41), .CLK(clk), .Q(
        decodedPacket3_o[38]) );
  DFFX1 \decodedPacket3_o_reg[37]  ( .D(n40), .CLK(clk), .Q(
        decodedPacket3_o[37]) );
  DFFX1 \decodedPacket3_o_reg[36]  ( .D(n39), .CLK(clk), .Q(
        decodedPacket3_o[36]) );
  DFFX1 \decodedPacket3_o_reg[35]  ( .D(n38), .CLK(clk), .Q(
        decodedPacket3_o[35]) );
  DFFX1 \decodedPacket3_o_reg[34]  ( .D(n37), .CLK(clk), .Q(
        decodedPacket3_o[34]) );
  DFFX1 \decodedPacket3_o_reg[33]  ( .D(n36), .CLK(clk), .Q(
        decodedPacket3_o[33]) );
  DFFX1 \decodedPacket3_o_reg[32]  ( .D(n35), .CLK(clk), .Q(
        decodedPacket3_o[32]) );
  DFFX1 \decodedPacket3_o_reg[31]  ( .D(n34), .CLK(clk), .Q(
        decodedPacket3_o[31]) );
  DFFX1 \decodedPacket3_o_reg[30]  ( .D(n33), .CLK(clk), .Q(
        decodedPacket3_o[30]) );
  DFFX1 \decodedPacket3_o_reg[29]  ( .D(n32), .CLK(clk), .Q(
        decodedPacket3_o[29]) );
  DFFX1 \decodedPacket3_o_reg[28]  ( .D(n31), .CLK(clk), .Q(
        decodedPacket3_o[28]) );
  DFFX1 \decodedPacket3_o_reg[27]  ( .D(n30), .CLK(clk), .Q(
        decodedPacket3_o[27]) );
  DFFX1 \decodedPacket3_o_reg[26]  ( .D(n29), .CLK(clk), .Q(
        decodedPacket3_o[26]) );
  DFFX1 \decodedPacket3_o_reg[25]  ( .D(n28), .CLK(clk), .Q(
        decodedPacket3_o[25]) );
  DFFX1 \decodedPacket3_o_reg[24]  ( .D(n27), .CLK(clk), .Q(
        decodedPacket3_o[24]) );
  DFFX1 \decodedPacket3_o_reg[23]  ( .D(n26), .CLK(clk), .Q(
        decodedPacket3_o[23]) );
  DFFX1 \decodedPacket3_o_reg[22]  ( .D(n25), .CLK(clk), .Q(
        decodedPacket3_o[22]) );
  DFFX1 \decodedPacket3_o_reg[21]  ( .D(n24), .CLK(clk), .Q(
        decodedPacket3_o[21]) );
  DFFX1 \decodedPacket3_o_reg[20]  ( .D(n23), .CLK(clk), .Q(
        decodedPacket3_o[20]) );
  DFFX1 \decodedPacket3_o_reg[19]  ( .D(n22), .CLK(clk), .Q(
        decodedPacket3_o[19]) );
  DFFX1 \decodedPacket3_o_reg[18]  ( .D(n21), .CLK(clk), .Q(
        decodedPacket3_o[18]) );
  DFFX1 \decodedPacket3_o_reg[17]  ( .D(n20), .CLK(clk), .Q(
        decodedPacket3_o[17]) );
  DFFX1 \decodedPacket3_o_reg[16]  ( .D(n19), .CLK(clk), .Q(
        decodedPacket3_o[16]) );
  DFFX1 \decodedPacket3_o_reg[15]  ( .D(n18), .CLK(clk), .Q(
        decodedPacket3_o[15]) );
  DFFX1 \decodedPacket3_o_reg[14]  ( .D(n17), .CLK(clk), .Q(
        decodedPacket3_o[14]) );
  DFFX1 \decodedPacket3_o_reg[13]  ( .D(n16), .CLK(clk), .Q(
        decodedPacket3_o[13]) );
  DFFX1 \decodedPacket3_o_reg[12]  ( .D(n15), .CLK(clk), .Q(
        decodedPacket3_o[12]) );
  DFFX1 \decodedPacket3_o_reg[11]  ( .D(n14), .CLK(clk), .Q(
        decodedPacket3_o[11]) );
  DFFX1 \decodedPacket3_o_reg[10]  ( .D(n13), .CLK(clk), .Q(
        decodedPacket3_o[10]) );
  DFFX1 \decodedPacket3_o_reg[9]  ( .D(n12), .CLK(clk), .Q(decodedPacket3_o[9]) );
  DFFX1 \decodedPacket3_o_reg[8]  ( .D(n11), .CLK(clk), .Q(decodedPacket3_o[8]) );
  DFFX1 \decodedPacket3_o_reg[7]  ( .D(n10), .CLK(clk), .Q(decodedPacket3_o[7]) );
  DFFX1 \decodedPacket3_o_reg[6]  ( .D(n9), .CLK(clk), .Q(decodedPacket3_o[6])
         );
  DFFX1 \decodedPacket3_o_reg[5]  ( .D(n8), .CLK(clk), .Q(decodedPacket3_o[5])
         );
  DFFX1 \decodedPacket3_o_reg[4]  ( .D(n7), .CLK(clk), .Q(decodedPacket3_o[4])
         );
  DFFX1 \decodedPacket3_o_reg[3]  ( .D(n6), .CLK(clk), .Q(decodedPacket3_o[3])
         );
  DFFX1 \decodedPacket3_o_reg[2]  ( .D(n5), .CLK(clk), .Q(decodedPacket3_o[2])
         );
  DFFX1 \decodedPacket3_o_reg[1]  ( .D(n4), .CLK(clk), .Q(decodedPacket3_o[1])
         );
  DFFX1 \decodedPacket3_o_reg[0]  ( .D(n3), .CLK(clk), .Q(decodedPacket3_o[0])
         );
  AO22X1 U2 ( .IN1(decodedPacket3_o[0]), .IN2(n577), .IN3(decodedPacket3_i[0]), 
        .IN4(n540), .Q(n3) );
  AO22X1 U3 ( .IN1(decodedPacket3_o[1]), .IN2(n577), .IN3(decodedPacket3_i[1]), 
        .IN4(n540), .Q(n4) );
  AO22X1 U4 ( .IN1(decodedPacket3_o[2]), .IN2(n577), .IN3(decodedPacket3_i[2]), 
        .IN4(n540), .Q(n5) );
  AO22X1 U5 ( .IN1(decodedPacket3_o[3]), .IN2(n577), .IN3(decodedPacket3_i[3]), 
        .IN4(n540), .Q(n6) );
  AO22X1 U6 ( .IN1(decodedPacket3_o[4]), .IN2(n576), .IN3(decodedPacket3_i[4]), 
        .IN4(n540), .Q(n7) );
  AO22X1 U7 ( .IN1(decodedPacket3_o[5]), .IN2(n576), .IN3(decodedPacket3_i[5]), 
        .IN4(n540), .Q(n8) );
  AO22X1 U8 ( .IN1(decodedPacket3_o[6]), .IN2(n576), .IN3(decodedPacket3_i[6]), 
        .IN4(n540), .Q(n9) );
  AO22X1 U9 ( .IN1(decodedPacket3_o[7]), .IN2(n576), .IN3(decodedPacket3_i[7]), 
        .IN4(n540), .Q(n10) );
  AO22X1 U10 ( .IN1(decodedPacket3_o[8]), .IN2(n576), .IN3(decodedPacket3_i[8]), .IN4(n540), .Q(n11) );
  AO22X1 U11 ( .IN1(decodedPacket3_o[9]), .IN2(n576), .IN3(decodedPacket3_i[9]), .IN4(n540), .Q(n12) );
  AO22X1 U12 ( .IN1(decodedPacket3_o[10]), .IN2(n576), .IN3(
        decodedPacket3_i[10]), .IN4(n540), .Q(n13) );
  AO22X1 U13 ( .IN1(decodedPacket3_o[11]), .IN2(n576), .IN3(
        decodedPacket3_i[11]), .IN4(n540), .Q(n14) );
  AO22X1 U14 ( .IN1(decodedPacket3_o[12]), .IN2(n576), .IN3(
        decodedPacket3_i[12]), .IN4(n540), .Q(n15) );
  AO22X1 U15 ( .IN1(decodedPacket3_o[13]), .IN2(n576), .IN3(
        decodedPacket3_i[13]), .IN4(n540), .Q(n16) );
  AO22X1 U16 ( .IN1(decodedPacket3_o[14]), .IN2(n576), .IN3(
        decodedPacket3_i[14]), .IN4(n540), .Q(n17) );
  AO22X1 U17 ( .IN1(decodedPacket3_o[15]), .IN2(n576), .IN3(
        decodedPacket3_i[15]), .IN4(n539), .Q(n18) );
  AO22X1 U18 ( .IN1(decodedPacket3_o[16]), .IN2(n568), .IN3(
        decodedPacket3_i[16]), .IN4(n539), .Q(n19) );
  AO22X1 U19 ( .IN1(decodedPacket3_o[17]), .IN2(n569), .IN3(
        decodedPacket3_i[17]), .IN4(n539), .Q(n20) );
  AO22X1 U20 ( .IN1(decodedPacket3_o[18]), .IN2(n570), .IN3(
        decodedPacket3_i[18]), .IN4(n539), .Q(n21) );
  AO22X1 U21 ( .IN1(decodedPacket3_o[19]), .IN2(n564), .IN3(
        decodedPacket3_i[19]), .IN4(n539), .Q(n22) );
  AO22X1 U22 ( .IN1(decodedPacket3_o[20]), .IN2(n565), .IN3(
        decodedPacket3_i[20]), .IN4(n539), .Q(n23) );
  AO22X1 U23 ( .IN1(decodedPacket3_o[21]), .IN2(n566), .IN3(
        decodedPacket3_i[21]), .IN4(n539), .Q(n24) );
  AO22X1 U24 ( .IN1(decodedPacket3_o[22]), .IN2(n567), .IN3(
        decodedPacket3_i[22]), .IN4(n539), .Q(n25) );
  AO22X1 U25 ( .IN1(decodedPacket3_o[23]), .IN2(n568), .IN3(
        decodedPacket3_i[23]), .IN4(n539), .Q(n26) );
  AO22X1 U26 ( .IN1(decodedPacket3_o[24]), .IN2(n569), .IN3(
        decodedPacket3_i[24]), .IN4(n539), .Q(n27) );
  AO22X1 U27 ( .IN1(decodedPacket3_o[25]), .IN2(n570), .IN3(
        decodedPacket3_i[25]), .IN4(n539), .Q(n28) );
  AO22X1 U28 ( .IN1(decodedPacket3_o[26]), .IN2(n563), .IN3(
        decodedPacket3_i[26]), .IN4(n539), .Q(n29) );
  AO22X1 U29 ( .IN1(decodedPacket3_o[27]), .IN2(n565), .IN3(
        decodedPacket3_i[27]), .IN4(n539), .Q(n30) );
  AO22X1 U30 ( .IN1(decodedPacket3_o[28]), .IN2(n575), .IN3(
        decodedPacket3_i[28]), .IN4(n539), .Q(n31) );
  AO22X1 U31 ( .IN1(decodedPacket3_o[29]), .IN2(n575), .IN3(
        decodedPacket3_i[29]), .IN4(n539), .Q(n32) );
  AO22X1 U32 ( .IN1(decodedPacket3_o[30]), .IN2(n575), .IN3(
        decodedPacket3_i[30]), .IN4(n539), .Q(n33) );
  AO22X1 U33 ( .IN1(decodedPacket3_o[31]), .IN2(n575), .IN3(
        decodedPacket3_i[31]), .IN4(n539), .Q(n34) );
  AO22X1 U34 ( .IN1(decodedPacket3_o[32]), .IN2(n575), .IN3(
        decodedPacket3_i[32]), .IN4(n539), .Q(n35) );
  AO22X1 U35 ( .IN1(decodedPacket3_o[33]), .IN2(n575), .IN3(
        decodedPacket3_i[33]), .IN4(n539), .Q(n36) );
  AO22X1 U36 ( .IN1(decodedPacket3_o[34]), .IN2(n575), .IN3(
        decodedPacket3_i[34]), .IN4(n538), .Q(n37) );
  AO22X1 U37 ( .IN1(decodedPacket3_o[35]), .IN2(n575), .IN3(
        decodedPacket3_i[35]), .IN4(n538), .Q(n38) );
  AO22X1 U38 ( .IN1(decodedPacket3_o[36]), .IN2(n575), .IN3(
        decodedPacket3_i[36]), .IN4(n538), .Q(n39) );
  AO22X1 U39 ( .IN1(decodedPacket3_o[37]), .IN2(n575), .IN3(
        decodedPacket3_i[37]), .IN4(n538), .Q(n40) );
  AO22X1 U40 ( .IN1(decodedPacket3_o[38]), .IN2(n575), .IN3(
        decodedPacket3_i[38]), .IN4(n538), .Q(n41) );
  AO22X1 U41 ( .IN1(decodedPacket3_o[39]), .IN2(n575), .IN3(
        decodedPacket3_i[39]), .IN4(n538), .Q(n42) );
  AO22X1 U42 ( .IN1(decodedPacket3_o[40]), .IN2(n547), .IN3(
        decodedPacket3_i[40]), .IN4(n538), .Q(n43) );
  AO22X1 U43 ( .IN1(decodedPacket3_o[41]), .IN2(n546), .IN3(
        decodedPacket3_i[41]), .IN4(n538), .Q(n44) );
  AO22X1 U44 ( .IN1(decodedPacket3_o[42]), .IN2(n545), .IN3(
        decodedPacket3_i[42]), .IN4(n538), .Q(n45) );
  AO22X1 U45 ( .IN1(decodedPacket3_o[43]), .IN2(n544), .IN3(
        decodedPacket3_i[43]), .IN4(n538), .Q(n46) );
  AO22X1 U46 ( .IN1(decodedPacket3_o[44]), .IN2(n543), .IN3(
        decodedPacket3_i[44]), .IN4(n538), .Q(n47) );
  AO22X1 U47 ( .IN1(decodedPacket3_o[45]), .IN2(n542), .IN3(
        decodedPacket3_i[45]), .IN4(n538), .Q(n48) );
  AO22X1 U48 ( .IN1(decodedPacket3_o[46]), .IN2(n541), .IN3(
        decodedPacket3_i[46]), .IN4(n538), .Q(n49) );
  AO22X1 U49 ( .IN1(decodedPacket3_o[47]), .IN2(n577), .IN3(
        decodedPacket3_i[47]), .IN4(n538), .Q(n50) );
  AO22X1 U50 ( .IN1(decodedPacket3_o[48]), .IN2(n580), .IN3(
        decodedPacket3_i[48]), .IN4(n538), .Q(n51) );
  AO22X1 U51 ( .IN1(decodedPacket3_o[49]), .IN2(n577), .IN3(
        decodedPacket3_i[49]), .IN4(n538), .Q(n52) );
  AO22X1 U52 ( .IN1(decodedPacket3_o[50]), .IN2(n577), .IN3(
        decodedPacket3_i[50]), .IN4(n538), .Q(n53) );
  AO22X1 U53 ( .IN1(decodedPacket3_o[51]), .IN2(n580), .IN3(
        decodedPacket3_i[51]), .IN4(n538), .Q(n54) );
  AO22X1 U54 ( .IN1(decodedPacket3_o[52]), .IN2(n574), .IN3(
        decodedPacket3_i[52]), .IN4(n538), .Q(n55) );
  AO22X1 U55 ( .IN1(decodedPacket3_o[53]), .IN2(n574), .IN3(
        decodedPacket3_i[53]), .IN4(n516), .Q(n56) );
  AO22X1 U56 ( .IN1(decodedPacket3_o[54]), .IN2(n574), .IN3(
        decodedPacket3_i[54]), .IN4(n516), .Q(n57) );
  AO22X1 U57 ( .IN1(decodedPacket3_o[55]), .IN2(n574), .IN3(
        decodedPacket3_i[55]), .IN4(n538), .Q(n58) );
  AO22X1 U58 ( .IN1(decodedPacket3_o[56]), .IN2(n574), .IN3(
        decodedPacket3_i[56]), .IN4(n539), .Q(n59) );
  AO22X1 U59 ( .IN1(decodedPacket3_o[57]), .IN2(n574), .IN3(
        decodedPacket3_i[57]), .IN4(n540), .Q(n60) );
  AO22X1 U60 ( .IN1(decodedPacket3_o[58]), .IN2(n574), .IN3(
        decodedPacket3_i[58]), .IN4(n511), .Q(n61) );
  AO22X1 U61 ( .IN1(decodedPacket3_o[59]), .IN2(n574), .IN3(
        decodedPacket3_i[59]), .IN4(n513), .Q(n62) );
  AO22X1 U62 ( .IN1(decodedPacket3_o[60]), .IN2(n574), .IN3(
        decodedPacket3_i[60]), .IN4(n527), .Q(n63) );
  AO22X1 U63 ( .IN1(decodedPacket3_o[61]), .IN2(n574), .IN3(
        decodedPacket3_i[61]), .IN4(n514), .Q(n64) );
  AO22X1 U64 ( .IN1(decodedPacket3_o[62]), .IN2(n574), .IN3(
        decodedPacket3_i[62]), .IN4(n517), .Q(n65) );
  AO22X1 U65 ( .IN1(decodedPacket3_o[63]), .IN2(n574), .IN3(
        decodedPacket3_i[63]), .IN4(n516), .Q(n66) );
  AO22X1 U66 ( .IN1(decodedPacket3_o[64]), .IN2(n573), .IN3(
        decodedPacket3_i[64]), .IN4(n516), .Q(n67) );
  AO22X1 U67 ( .IN1(decodedPacket3_o[65]), .IN2(n573), .IN3(
        decodedPacket3_i[65]), .IN4(n511), .Q(n68) );
  AO22X1 U68 ( .IN1(decodedPacket3_o[66]), .IN2(n573), .IN3(
        decodedPacket3_i[66]), .IN4(n513), .Q(n69) );
  AO22X1 U69 ( .IN1(decodedPacket3_o[67]), .IN2(n573), .IN3(
        decodedPacket3_i[67]), .IN4(n528), .Q(n70) );
  AO22X1 U70 ( .IN1(decodedPacket3_o[68]), .IN2(n573), .IN3(
        decodedPacket3_i[68]), .IN4(n535), .Q(n71) );
  AO22X1 U71 ( .IN1(decodedPacket3_o[69]), .IN2(n573), .IN3(
        decodedPacket3_i[69]), .IN4(n530), .Q(n72) );
  AO22X1 U72 ( .IN1(decodedPacket3_o[70]), .IN2(n573), .IN3(
        decodedPacket3_i[70]), .IN4(n521), .Q(n73) );
  AO22X1 U73 ( .IN1(decodedPacket3_o[71]), .IN2(n573), .IN3(
        decodedPacket3_i[71]), .IN4(n522), .Q(n74) );
  AO22X1 U74 ( .IN1(decodedPacket3_o[72]), .IN2(n573), .IN3(
        decodedPacket3_i[72]), .IN4(n537), .Q(n75) );
  AO22X1 U75 ( .IN1(decodedPacket3_o[73]), .IN2(n573), .IN3(
        decodedPacket3_i[73]), .IN4(n537), .Q(n76) );
  AO22X1 U76 ( .IN1(decodedPacket3_o[74]), .IN2(n573), .IN3(
        decodedPacket3_i[74]), .IN4(n537), .Q(n77) );
  AO22X1 U77 ( .IN1(decodedPacket3_o[75]), .IN2(n573), .IN3(
        decodedPacket3_i[75]), .IN4(n537), .Q(n78) );
  AO22X1 U78 ( .IN1(decodedPacket3_o[76]), .IN2(n577), .IN3(
        decodedPacket3_i[76]), .IN4(n537), .Q(n79) );
  AO22X1 U79 ( .IN1(decodedPacket3_o[77]), .IN2(n577), .IN3(
        decodedPacket3_i[77]), .IN4(n537), .Q(n80) );
  AO22X1 U80 ( .IN1(decodedPacket3_o[78]), .IN2(n577), .IN3(
        decodedPacket3_i[78]), .IN4(n537), .Q(n81) );
  AO22X1 U81 ( .IN1(decodedPacket3_o[79]), .IN2(n577), .IN3(
        decodedPacket3_i[79]), .IN4(n537), .Q(n82) );
  AO22X1 U82 ( .IN1(decodedPacket3_o[80]), .IN2(n547), .IN3(
        decodedPacket3_i[80]), .IN4(n537), .Q(n83) );
  AO22X1 U83 ( .IN1(decodedPacket3_o[81]), .IN2(n546), .IN3(
        decodedPacket3_i[81]), .IN4(n537), .Q(n84) );
  AO22X1 U84 ( .IN1(decodedPacket3_o[82]), .IN2(n545), .IN3(
        decodedPacket3_i[82]), .IN4(n537), .Q(n85) );
  AO22X1 U85 ( .IN1(decodedPacket3_o[83]), .IN2(n544), .IN3(
        decodedPacket3_i[83]), .IN4(n537), .Q(n86) );
  AO22X1 U86 ( .IN1(decodedPacket3_o[84]), .IN2(n543), .IN3(
        decodedPacket3_i[84]), .IN4(n537), .Q(n87) );
  AO22X1 U87 ( .IN1(decodedPacket3_o[85]), .IN2(n542), .IN3(
        decodedPacket3_i[85]), .IN4(n537), .Q(n88) );
  AO22X1 U88 ( .IN1(decodedPacket3_o[86]), .IN2(n541), .IN3(
        decodedPacket3_i[86]), .IN4(n537), .Q(n89) );
  AO22X1 U89 ( .IN1(decodedPacket3_o[87]), .IN2(n577), .IN3(
        decodedPacket3_i[87]), .IN4(n537), .Q(n90) );
  AO22X1 U90 ( .IN1(decodedPacket3_o[88]), .IN2(n577), .IN3(
        decodedPacket3_i[88]), .IN4(n537), .Q(n91) );
  AO22X1 U91 ( .IN1(decodedPacket3_o[89]), .IN2(n572), .IN3(
        decodedPacket3_i[89]), .IN4(n537), .Q(n92) );
  AO22X1 U92 ( .IN1(decodedPacket3_o[90]), .IN2(n571), .IN3(
        decodedPacket3_i[90]), .IN4(n537), .Q(n93) );
  AO22X1 U93 ( .IN1(decodedPacket3_o[91]), .IN2(n573), .IN3(
        decodedPacket3_i[91]), .IN4(n536), .Q(n94) );
  AO22X1 U94 ( .IN1(decodedPacket3_o[92]), .IN2(n575), .IN3(
        decodedPacket3_i[92]), .IN4(n536), .Q(n95) );
  AO22X1 U95 ( .IN1(decodedPacket3_o[93]), .IN2(n574), .IN3(
        decodedPacket3_i[93]), .IN4(n536), .Q(n96) );
  AO22X1 U96 ( .IN1(decodedPacket3_o[94]), .IN2(n577), .IN3(
        decodedPacket3_i[94]), .IN4(n536), .Q(n97) );
  AO22X1 U97 ( .IN1(decodedPacket3_o[95]), .IN2(n576), .IN3(
        decodedPacket3_i[95]), .IN4(n536), .Q(n98) );
  AO22X1 U98 ( .IN1(decodedPacket3_o[96]), .IN2(n567), .IN3(
        decodedPacket3_i[96]), .IN4(n536), .Q(n99) );
  AO22X1 U99 ( .IN1(decodedPacket3_o[97]), .IN2(n578), .IN3(
        decodedPacket3_i[97]), .IN4(n536), .Q(n100) );
  AO22X1 U100 ( .IN1(decodedPacket3_o[98]), .IN2(n547), .IN3(
        decodedPacket3_i[98]), .IN4(n536), .Q(n101) );
  AO22X1 U101 ( .IN1(decodedPacket3_o[99]), .IN2(n546), .IN3(
        decodedPacket3_i[99]), .IN4(n536), .Q(n102) );
  AO22X1 U102 ( .IN1(decodedPacket3_o[100]), .IN2(n572), .IN3(
        decodedPacket3_i[100]), .IN4(n536), .Q(n103) );
  AO22X1 U103 ( .IN1(decodedPacket3_o[101]), .IN2(n571), .IN3(
        decodedPacket3_i[101]), .IN4(n536), .Q(n104) );
  AO22X1 U104 ( .IN1(decodedPacket3_o[102]), .IN2(n573), .IN3(
        decodedPacket3_i[102]), .IN4(n536), .Q(n105) );
  AO22X1 U105 ( .IN1(decodedPacket3_o[103]), .IN2(n576), .IN3(
        decodedPacket3_i[103]), .IN4(n536), .Q(n106) );
  AO22X1 U106 ( .IN1(decodedPacket3_o[104]), .IN2(n566), .IN3(
        decodedPacket3_i[104]), .IN4(n536), .Q(n107) );
  AO22X1 U107 ( .IN1(decodedPacket3_o[105]), .IN2(n575), .IN3(
        decodedPacket3_i[105]), .IN4(n536), .Q(n108) );
  AO22X1 U108 ( .IN1(decodedPacket3_o[106]), .IN2(n574), .IN3(
        decodedPacket3_i[106]), .IN4(n536), .Q(n109) );
  AO22X1 U109 ( .IN1(decodedPacket3_o[107]), .IN2(n578), .IN3(
        decodedPacket3_i[107]), .IN4(n536), .Q(n110) );
  AO22X1 U110 ( .IN1(decodedPacket3_o[108]), .IN2(n545), .IN3(
        decodedPacket3_i[108]), .IN4(n536), .Q(n111) );
  AO22X1 U111 ( .IN1(decodedPacket3_o[109]), .IN2(n544), .IN3(
        decodedPacket3_i[109]), .IN4(n536), .Q(n112) );
  AO22X1 U112 ( .IN1(decodedPacket3_o[110]), .IN2(n543), .IN3(
        decodedPacket3_i[110]), .IN4(n535), .Q(n113) );
  AO22X1 U113 ( .IN1(decodedPacket3_o[111]), .IN2(n542), .IN3(
        decodedPacket3_i[111]), .IN4(n535), .Q(n114) );
  AO22X1 U114 ( .IN1(decodedPacket3_o[112]), .IN2(n572), .IN3(
        decodedPacket3_i[112]), .IN4(n535), .Q(n115) );
  AO22X1 U115 ( .IN1(decodedPacket3_o[113]), .IN2(n572), .IN3(
        decodedPacket3_i[113]), .IN4(n535), .Q(n116) );
  AO22X1 U116 ( .IN1(decodedPacket3_o[114]), .IN2(n572), .IN3(
        decodedPacket3_i[114]), .IN4(n535), .Q(n117) );
  AO22X1 U117 ( .IN1(decodedPacket3_o[115]), .IN2(n572), .IN3(
        decodedPacket3_i[115]), .IN4(n535), .Q(n118) );
  AO22X1 U118 ( .IN1(decodedPacket3_o[116]), .IN2(n572), .IN3(
        decodedPacket3_i[116]), .IN4(n535), .Q(n119) );
  AO22X1 U119 ( .IN1(decodedPacket3_o[117]), .IN2(n572), .IN3(
        decodedPacket3_i[117]), .IN4(n535), .Q(n120) );
  AO22X1 U120 ( .IN1(decodedPacket3_o[118]), .IN2(n572), .IN3(
        decodedPacket3_i[118]), .IN4(n535), .Q(n121) );
  AO22X1 U121 ( .IN1(decodedPacket3_o[119]), .IN2(n572), .IN3(
        decodedPacket3_i[119]), .IN4(n535), .Q(n122) );
  AO22X1 U122 ( .IN1(decodedPacket3_o[120]), .IN2(n572), .IN3(
        decodedPacket3_i[120]), .IN4(n535), .Q(n123) );
  AO22X1 U123 ( .IN1(decodedPacket3_o[121]), .IN2(n572), .IN3(
        decodedPacket3_i[121]), .IN4(n535), .Q(n124) );
  AO22X1 U124 ( .IN1(decodedPacket3_o[122]), .IN2(n572), .IN3(
        decodedPacket3_i[122]), .IN4(n535), .Q(n125) );
  AO22X1 U125 ( .IN1(decodedPacket3_o[123]), .IN2(n572), .IN3(
        decodedPacket3_i[123]), .IN4(n535), .Q(n126) );
  AO22X1 U126 ( .IN1(decodedPacket3_o[124]), .IN2(n571), .IN3(
        decodedPacket3_i[124]), .IN4(n535), .Q(n127) );
  AO22X1 U127 ( .IN1(decodedPacket3_o[125]), .IN2(n571), .IN3(
        decodedPacket3_i[125]), .IN4(n535), .Q(n128) );
  AO22X1 U128 ( .IN1(decodedPacket2_o[0]), .IN2(n571), .IN3(
        decodedPacket2_i[0]), .IN4(n535), .Q(n129) );
  AO22X1 U129 ( .IN1(decodedPacket2_o[1]), .IN2(n571), .IN3(
        decodedPacket2_i[1]), .IN4(n535), .Q(n130) );
  AO22X1 U130 ( .IN1(decodedPacket2_o[2]), .IN2(n571), .IN3(
        decodedPacket2_i[2]), .IN4(n535), .Q(n131) );
  AO22X1 U131 ( .IN1(decodedPacket2_o[3]), .IN2(n571), .IN3(
        decodedPacket2_i[3]), .IN4(n534), .Q(n132) );
  AO22X1 U132 ( .IN1(decodedPacket2_o[4]), .IN2(n571), .IN3(
        decodedPacket2_i[4]), .IN4(n534), .Q(n133) );
  AO22X1 U133 ( .IN1(decodedPacket2_o[5]), .IN2(n571), .IN3(
        decodedPacket2_i[5]), .IN4(n534), .Q(n134) );
  AO22X1 U134 ( .IN1(decodedPacket2_o[6]), .IN2(n571), .IN3(
        decodedPacket2_i[6]), .IN4(n534), .Q(n135) );
  AO22X1 U135 ( .IN1(decodedPacket2_o[7]), .IN2(n571), .IN3(
        decodedPacket2_i[7]), .IN4(n534), .Q(n136) );
  AO22X1 U136 ( .IN1(decodedPacket2_o[8]), .IN2(n571), .IN3(
        decodedPacket2_i[8]), .IN4(n534), .Q(n137) );
  AO22X1 U137 ( .IN1(decodedPacket2_o[9]), .IN2(n571), .IN3(
        decodedPacket2_i[9]), .IN4(n534), .Q(n138) );
  AO22X1 U138 ( .IN1(decodedPacket2_o[10]), .IN2(n570), .IN3(
        decodedPacket2_i[10]), .IN4(n534), .Q(n139) );
  AO22X1 U139 ( .IN1(decodedPacket2_o[11]), .IN2(n570), .IN3(
        decodedPacket2_i[11]), .IN4(n534), .Q(n140) );
  AO22X1 U140 ( .IN1(decodedPacket2_o[12]), .IN2(n570), .IN3(
        decodedPacket2_i[12]), .IN4(n534), .Q(n141) );
  AO22X1 U141 ( .IN1(decodedPacket2_o[13]), .IN2(n570), .IN3(
        decodedPacket2_i[13]), .IN4(n534), .Q(n142) );
  AO22X1 U142 ( .IN1(decodedPacket2_o[14]), .IN2(n570), .IN3(
        decodedPacket2_i[14]), .IN4(n534), .Q(n143) );
  AO22X1 U143 ( .IN1(decodedPacket2_o[15]), .IN2(n570), .IN3(
        decodedPacket2_i[15]), .IN4(n534), .Q(n144) );
  AO22X1 U144 ( .IN1(decodedPacket2_o[16]), .IN2(n570), .IN3(
        decodedPacket2_i[16]), .IN4(n534), .Q(n145) );
  AO22X1 U145 ( .IN1(decodedPacket2_o[17]), .IN2(n570), .IN3(
        decodedPacket2_i[17]), .IN4(n534), .Q(n146) );
  AO22X1 U146 ( .IN1(decodedPacket2_o[18]), .IN2(n570), .IN3(
        decodedPacket2_i[18]), .IN4(n534), .Q(n147) );
  AO22X1 U147 ( .IN1(decodedPacket2_o[19]), .IN2(n570), .IN3(
        decodedPacket2_i[19]), .IN4(n534), .Q(n148) );
  AO22X1 U148 ( .IN1(decodedPacket2_o[20]), .IN2(n570), .IN3(
        decodedPacket2_i[20]), .IN4(n534), .Q(n149) );
  AO22X1 U149 ( .IN1(decodedPacket2_o[21]), .IN2(n570), .IN3(
        decodedPacket2_i[21]), .IN4(n534), .Q(n150) );
  AO22X1 U150 ( .IN1(decodedPacket2_o[22]), .IN2(n569), .IN3(
        decodedPacket2_i[22]), .IN4(n533), .Q(n151) );
  AO22X1 U151 ( .IN1(decodedPacket2_o[23]), .IN2(n569), .IN3(
        decodedPacket2_i[23]), .IN4(n533), .Q(n152) );
  AO22X1 U152 ( .IN1(decodedPacket2_o[24]), .IN2(n569), .IN3(
        decodedPacket2_i[24]), .IN4(n533), .Q(n153) );
  AO22X1 U153 ( .IN1(decodedPacket2_o[25]), .IN2(n569), .IN3(
        decodedPacket2_i[25]), .IN4(n533), .Q(n154) );
  AO22X1 U154 ( .IN1(decodedPacket2_o[26]), .IN2(n569), .IN3(
        decodedPacket2_i[26]), .IN4(n533), .Q(n155) );
  AO22X1 U155 ( .IN1(decodedPacket2_o[27]), .IN2(n569), .IN3(
        decodedPacket2_i[27]), .IN4(n533), .Q(n156) );
  AO22X1 U156 ( .IN1(decodedPacket2_o[28]), .IN2(n569), .IN3(
        decodedPacket2_i[28]), .IN4(n533), .Q(n157) );
  AO22X1 U157 ( .IN1(decodedPacket2_o[29]), .IN2(n569), .IN3(
        decodedPacket2_i[29]), .IN4(n533), .Q(n158) );
  AO22X1 U158 ( .IN1(decodedPacket2_o[30]), .IN2(n569), .IN3(
        decodedPacket2_i[30]), .IN4(n533), .Q(n159) );
  AO22X1 U159 ( .IN1(decodedPacket2_o[31]), .IN2(n569), .IN3(
        decodedPacket2_i[31]), .IN4(n533), .Q(n160) );
  AO22X1 U160 ( .IN1(decodedPacket2_o[32]), .IN2(n569), .IN3(
        decodedPacket2_i[32]), .IN4(n533), .Q(n161) );
  AO22X1 U161 ( .IN1(decodedPacket2_o[33]), .IN2(n569), .IN3(
        decodedPacket2_i[33]), .IN4(n533), .Q(n162) );
  AO22X1 U162 ( .IN1(decodedPacket2_o[34]), .IN2(n568), .IN3(
        decodedPacket2_i[34]), .IN4(n533), .Q(n163) );
  AO22X1 U163 ( .IN1(decodedPacket2_o[35]), .IN2(n568), .IN3(
        decodedPacket2_i[35]), .IN4(n533), .Q(n164) );
  AO22X1 U164 ( .IN1(decodedPacket2_o[36]), .IN2(n568), .IN3(
        decodedPacket2_i[36]), .IN4(n533), .Q(n165) );
  AO22X1 U165 ( .IN1(decodedPacket2_o[37]), .IN2(n568), .IN3(
        decodedPacket2_i[37]), .IN4(n533), .Q(n166) );
  AO22X1 U166 ( .IN1(decodedPacket2_o[38]), .IN2(n568), .IN3(
        decodedPacket2_i[38]), .IN4(n533), .Q(n167) );
  AO22X1 U167 ( .IN1(decodedPacket2_o[39]), .IN2(n568), .IN3(
        decodedPacket2_i[39]), .IN4(n533), .Q(n168) );
  AO22X1 U168 ( .IN1(decodedPacket2_o[40]), .IN2(n568), .IN3(
        decodedPacket2_i[40]), .IN4(n533), .Q(n169) );
  AO22X1 U169 ( .IN1(decodedPacket2_o[41]), .IN2(n568), .IN3(
        decodedPacket2_i[41]), .IN4(n532), .Q(n170) );
  AO22X1 U170 ( .IN1(decodedPacket2_o[42]), .IN2(n568), .IN3(
        decodedPacket2_i[42]), .IN4(n532), .Q(n171) );
  AO22X1 U171 ( .IN1(decodedPacket2_o[43]), .IN2(n568), .IN3(
        decodedPacket2_i[43]), .IN4(n532), .Q(n172) );
  AO22X1 U172 ( .IN1(decodedPacket2_o[44]), .IN2(n568), .IN3(
        decodedPacket2_i[44]), .IN4(n532), .Q(n173) );
  AO22X1 U173 ( .IN1(decodedPacket2_o[45]), .IN2(n568), .IN3(
        decodedPacket2_i[45]), .IN4(n532), .Q(n174) );
  AO22X1 U174 ( .IN1(decodedPacket2_o[46]), .IN2(n567), .IN3(
        decodedPacket2_i[46]), .IN4(n532), .Q(n175) );
  AO22X1 U175 ( .IN1(decodedPacket2_o[47]), .IN2(n567), .IN3(
        decodedPacket2_i[47]), .IN4(n532), .Q(n176) );
  AO22X1 U176 ( .IN1(decodedPacket2_o[48]), .IN2(n567), .IN3(
        decodedPacket2_i[48]), .IN4(n532), .Q(n177) );
  AO22X1 U177 ( .IN1(decodedPacket2_o[49]), .IN2(n567), .IN3(
        decodedPacket2_i[49]), .IN4(n532), .Q(n178) );
  AO22X1 U178 ( .IN1(decodedPacket2_o[50]), .IN2(n567), .IN3(
        decodedPacket2_i[50]), .IN4(n532), .Q(n179) );
  AO22X1 U179 ( .IN1(decodedPacket2_o[51]), .IN2(n567), .IN3(
        decodedPacket2_i[51]), .IN4(n532), .Q(n180) );
  AO22X1 U180 ( .IN1(decodedPacket2_o[52]), .IN2(n567), .IN3(
        decodedPacket2_i[52]), .IN4(n532), .Q(n181) );
  AO22X1 U181 ( .IN1(decodedPacket2_o[53]), .IN2(n567), .IN3(
        decodedPacket2_i[53]), .IN4(n532), .Q(n182) );
  AO22X1 U182 ( .IN1(decodedPacket2_o[54]), .IN2(n567), .IN3(
        decodedPacket2_i[54]), .IN4(n532), .Q(n183) );
  AO22X1 U183 ( .IN1(decodedPacket2_o[55]), .IN2(n567), .IN3(
        decodedPacket2_i[55]), .IN4(n532), .Q(n184) );
  AO22X1 U184 ( .IN1(decodedPacket2_o[56]), .IN2(n567), .IN3(
        decodedPacket2_i[56]), .IN4(n532), .Q(n185) );
  AO22X1 U185 ( .IN1(decodedPacket2_o[57]), .IN2(n567), .IN3(
        decodedPacket2_i[57]), .IN4(n532), .Q(n186) );
  AO22X1 U186 ( .IN1(decodedPacket2_o[58]), .IN2(n566), .IN3(
        decodedPacket2_i[58]), .IN4(n532), .Q(n187) );
  AO22X1 U187 ( .IN1(decodedPacket2_o[59]), .IN2(n566), .IN3(
        decodedPacket2_i[59]), .IN4(n532), .Q(n188) );
  AO22X1 U188 ( .IN1(decodedPacket2_o[60]), .IN2(n566), .IN3(
        decodedPacket2_i[60]), .IN4(n531), .Q(n189) );
  AO22X1 U189 ( .IN1(decodedPacket2_o[61]), .IN2(n566), .IN3(
        decodedPacket2_i[61]), .IN4(n531), .Q(n190) );
  AO22X1 U190 ( .IN1(decodedPacket2_o[62]), .IN2(n566), .IN3(
        decodedPacket2_i[62]), .IN4(n531), .Q(n191) );
  AO22X1 U191 ( .IN1(decodedPacket2_o[63]), .IN2(n566), .IN3(
        decodedPacket2_i[63]), .IN4(n531), .Q(n192) );
  AO22X1 U192 ( .IN1(decodedPacket2_o[64]), .IN2(n566), .IN3(
        decodedPacket2_i[64]), .IN4(n531), .Q(n193) );
  AO22X1 U193 ( .IN1(decodedPacket2_o[65]), .IN2(n566), .IN3(
        decodedPacket2_i[65]), .IN4(n531), .Q(n194) );
  AO22X1 U194 ( .IN1(decodedPacket2_o[66]), .IN2(n566), .IN3(
        decodedPacket2_i[66]), .IN4(n531), .Q(n195) );
  AO22X1 U195 ( .IN1(decodedPacket2_o[67]), .IN2(n566), .IN3(
        decodedPacket2_i[67]), .IN4(n531), .Q(n196) );
  AO22X1 U196 ( .IN1(decodedPacket2_o[68]), .IN2(n566), .IN3(
        decodedPacket2_i[68]), .IN4(n531), .Q(n197) );
  AO22X1 U197 ( .IN1(decodedPacket2_o[69]), .IN2(n566), .IN3(
        decodedPacket2_i[69]), .IN4(n531), .Q(n198) );
  AO22X1 U198 ( .IN1(decodedPacket2_o[70]), .IN2(n565), .IN3(
        decodedPacket2_i[70]), .IN4(n531), .Q(n199) );
  AO22X1 U199 ( .IN1(decodedPacket2_o[71]), .IN2(n565), .IN3(
        decodedPacket2_i[71]), .IN4(n531), .Q(n200) );
  AO22X1 U200 ( .IN1(decodedPacket2_o[72]), .IN2(n565), .IN3(
        decodedPacket2_i[72]), .IN4(n531), .Q(n201) );
  AO22X1 U201 ( .IN1(decodedPacket2_o[73]), .IN2(n565), .IN3(
        decodedPacket2_i[73]), .IN4(n531), .Q(n202) );
  AO22X1 U202 ( .IN1(decodedPacket2_o[74]), .IN2(n565), .IN3(
        decodedPacket2_i[74]), .IN4(n531), .Q(n203) );
  AO22X1 U203 ( .IN1(decodedPacket2_o[75]), .IN2(n565), .IN3(
        decodedPacket2_i[75]), .IN4(n531), .Q(n204) );
  AO22X1 U204 ( .IN1(decodedPacket2_o[76]), .IN2(n565), .IN3(
        decodedPacket2_i[76]), .IN4(n531), .Q(n205) );
  AO22X1 U205 ( .IN1(decodedPacket2_o[77]), .IN2(n565), .IN3(
        decodedPacket2_i[77]), .IN4(n531), .Q(n206) );
  AO22X1 U206 ( .IN1(decodedPacket2_o[78]), .IN2(n565), .IN3(
        decodedPacket2_i[78]), .IN4(n531), .Q(n207) );
  AO22X1 U207 ( .IN1(decodedPacket2_o[79]), .IN2(n565), .IN3(
        decodedPacket2_i[79]), .IN4(n530), .Q(n208) );
  AO22X1 U208 ( .IN1(decodedPacket2_o[80]), .IN2(n565), .IN3(
        decodedPacket2_i[80]), .IN4(n530), .Q(n209) );
  AO22X1 U209 ( .IN1(decodedPacket2_o[81]), .IN2(n565), .IN3(
        decodedPacket2_i[81]), .IN4(n530), .Q(n210) );
  AO22X1 U210 ( .IN1(decodedPacket2_o[82]), .IN2(n564), .IN3(
        decodedPacket2_i[82]), .IN4(n530), .Q(n211) );
  AO22X1 U211 ( .IN1(decodedPacket2_o[83]), .IN2(n564), .IN3(
        decodedPacket2_i[83]), .IN4(n530), .Q(n212) );
  AO22X1 U212 ( .IN1(decodedPacket2_o[84]), .IN2(n564), .IN3(
        decodedPacket2_i[84]), .IN4(n530), .Q(n213) );
  AO22X1 U213 ( .IN1(decodedPacket2_o[85]), .IN2(n564), .IN3(
        decodedPacket2_i[85]), .IN4(n530), .Q(n214) );
  AO22X1 U214 ( .IN1(decodedPacket2_o[86]), .IN2(n564), .IN3(
        decodedPacket2_i[86]), .IN4(n530), .Q(n215) );
  AO22X1 U215 ( .IN1(decodedPacket2_o[87]), .IN2(n564), .IN3(
        decodedPacket2_i[87]), .IN4(n530), .Q(n216) );
  AO22X1 U216 ( .IN1(decodedPacket2_o[88]), .IN2(n564), .IN3(
        decodedPacket2_i[88]), .IN4(n530), .Q(n217) );
  AO22X1 U217 ( .IN1(decodedPacket2_o[89]), .IN2(n564), .IN3(
        decodedPacket2_i[89]), .IN4(n530), .Q(n218) );
  AO22X1 U218 ( .IN1(decodedPacket2_o[90]), .IN2(n564), .IN3(
        decodedPacket2_i[90]), .IN4(n530), .Q(n219) );
  AO22X1 U219 ( .IN1(decodedPacket2_o[91]), .IN2(n564), .IN3(
        decodedPacket2_i[91]), .IN4(n530), .Q(n220) );
  AO22X1 U220 ( .IN1(decodedPacket2_o[92]), .IN2(n564), .IN3(
        decodedPacket2_i[92]), .IN4(n530), .Q(n221) );
  AO22X1 U221 ( .IN1(decodedPacket2_o[93]), .IN2(n564), .IN3(
        decodedPacket2_i[93]), .IN4(n530), .Q(n222) );
  AO22X1 U222 ( .IN1(decodedPacket2_o[94]), .IN2(n563), .IN3(
        decodedPacket2_i[94]), .IN4(n530), .Q(n223) );
  AO22X1 U223 ( .IN1(decodedPacket2_o[95]), .IN2(n563), .IN3(
        decodedPacket2_i[95]), .IN4(n530), .Q(n224) );
  AO22X1 U224 ( .IN1(decodedPacket2_o[96]), .IN2(n563), .IN3(
        decodedPacket2_i[96]), .IN4(n530), .Q(n225) );
  AO22X1 U225 ( .IN1(decodedPacket2_o[97]), .IN2(n563), .IN3(
        decodedPacket2_i[97]), .IN4(n530), .Q(n226) );
  AO22X1 U226 ( .IN1(decodedPacket2_o[98]), .IN2(n563), .IN3(
        decodedPacket2_i[98]), .IN4(n529), .Q(n227) );
  AO22X1 U227 ( .IN1(decodedPacket2_o[99]), .IN2(n563), .IN3(
        decodedPacket2_i[99]), .IN4(n529), .Q(n228) );
  AO22X1 U228 ( .IN1(decodedPacket2_o[100]), .IN2(n563), .IN3(
        decodedPacket2_i[100]), .IN4(n529), .Q(n229) );
  AO22X1 U229 ( .IN1(decodedPacket2_o[101]), .IN2(n563), .IN3(
        decodedPacket2_i[101]), .IN4(n529), .Q(n230) );
  AO22X1 U230 ( .IN1(decodedPacket2_o[102]), .IN2(n563), .IN3(
        decodedPacket2_i[102]), .IN4(n529), .Q(n231) );
  AO22X1 U231 ( .IN1(decodedPacket2_o[103]), .IN2(n563), .IN3(
        decodedPacket2_i[103]), .IN4(n529), .Q(n232) );
  AO22X1 U232 ( .IN1(decodedPacket2_o[104]), .IN2(n563), .IN3(
        decodedPacket2_i[104]), .IN4(n529), .Q(n233) );
  AO22X1 U233 ( .IN1(decodedPacket2_o[105]), .IN2(n563), .IN3(
        decodedPacket2_i[105]), .IN4(n529), .Q(n234) );
  AO22X1 U234 ( .IN1(decodedPacket2_o[106]), .IN2(n563), .IN3(
        decodedPacket2_i[106]), .IN4(n529), .Q(n235) );
  AO22X1 U235 ( .IN1(decodedPacket2_o[107]), .IN2(n564), .IN3(
        decodedPacket2_i[107]), .IN4(n529), .Q(n236) );
  AO22X1 U236 ( .IN1(decodedPacket2_o[108]), .IN2(n566), .IN3(
        decodedPacket2_i[108]), .IN4(n529), .Q(n237) );
  AO22X1 U237 ( .IN1(decodedPacket2_o[109]), .IN2(n567), .IN3(
        decodedPacket2_i[109]), .IN4(n529), .Q(n238) );
  AO22X1 U238 ( .IN1(decodedPacket2_o[110]), .IN2(n568), .IN3(
        decodedPacket2_i[110]), .IN4(n529), .Q(n239) );
  AO22X1 U239 ( .IN1(decodedPacket2_o[111]), .IN2(n569), .IN3(
        decodedPacket2_i[111]), .IN4(n529), .Q(n240) );
  AO22X1 U240 ( .IN1(decodedPacket2_o[112]), .IN2(n570), .IN3(
        decodedPacket2_i[112]), .IN4(n529), .Q(n241) );
  AO22X1 U241 ( .IN1(decodedPacket2_o[113]), .IN2(n565), .IN3(
        decodedPacket2_i[113]), .IN4(n529), .Q(n242) );
  AO22X1 U242 ( .IN1(decodedPacket2_o[114]), .IN2(n563), .IN3(
        decodedPacket2_i[114]), .IN4(n529), .Q(n243) );
  AO22X1 U243 ( .IN1(decodedPacket2_o[115]), .IN2(n564), .IN3(
        decodedPacket2_i[115]), .IN4(n529), .Q(n244) );
  AO22X1 U244 ( .IN1(decodedPacket2_o[116]), .IN2(n566), .IN3(
        decodedPacket2_i[116]), .IN4(n529), .Q(n245) );
  AO22X1 U245 ( .IN1(decodedPacket2_o[117]), .IN2(n567), .IN3(
        decodedPacket2_i[117]), .IN4(n528), .Q(n246) );
  AO22X1 U246 ( .IN1(decodedPacket2_o[118]), .IN2(n562), .IN3(
        decodedPacket2_i[118]), .IN4(n528), .Q(n247) );
  AO22X1 U247 ( .IN1(decodedPacket2_o[119]), .IN2(n562), .IN3(
        decodedPacket2_i[119]), .IN4(n528), .Q(n248) );
  AO22X1 U248 ( .IN1(decodedPacket2_o[120]), .IN2(n562), .IN3(
        decodedPacket2_i[120]), .IN4(n528), .Q(n249) );
  AO22X1 U249 ( .IN1(decodedPacket2_o[121]), .IN2(n562), .IN3(
        decodedPacket2_i[121]), .IN4(n528), .Q(n250) );
  AO22X1 U250 ( .IN1(decodedPacket2_o[122]), .IN2(n562), .IN3(
        decodedPacket2_i[122]), .IN4(n528), .Q(n251) );
  AO22X1 U251 ( .IN1(decodedPacket2_o[123]), .IN2(n562), .IN3(
        decodedPacket2_i[123]), .IN4(n528), .Q(n252) );
  AO22X1 U252 ( .IN1(decodedPacket2_o[124]), .IN2(n562), .IN3(
        decodedPacket2_i[124]), .IN4(n528), .Q(n253) );
  AO22X1 U253 ( .IN1(decodedPacket2_o[125]), .IN2(n562), .IN3(
        decodedPacket2_i[125]), .IN4(n528), .Q(n254) );
  AO22X1 U254 ( .IN1(decodedPacket1_o[0]), .IN2(n562), .IN3(
        decodedPacket1_i[0]), .IN4(n528), .Q(n255) );
  AO22X1 U255 ( .IN1(decodedPacket1_o[1]), .IN2(n562), .IN3(
        decodedPacket1_i[1]), .IN4(n528), .Q(n256) );
  AO22X1 U256 ( .IN1(decodedPacket1_o[2]), .IN2(n562), .IN3(
        decodedPacket1_i[2]), .IN4(n528), .Q(n257) );
  AO22X1 U257 ( .IN1(decodedPacket1_o[3]), .IN2(n562), .IN3(
        decodedPacket1_i[3]), .IN4(n528), .Q(n258) );
  AO22X1 U258 ( .IN1(decodedPacket1_o[4]), .IN2(n561), .IN3(
        decodedPacket1_i[4]), .IN4(n528), .Q(n259) );
  AO22X1 U259 ( .IN1(decodedPacket1_o[5]), .IN2(n561), .IN3(
        decodedPacket1_i[5]), .IN4(n528), .Q(n260) );
  AO22X1 U260 ( .IN1(decodedPacket1_o[6]), .IN2(n561), .IN3(
        decodedPacket1_i[6]), .IN4(n528), .Q(n261) );
  AO22X1 U261 ( .IN1(decodedPacket1_o[7]), .IN2(n561), .IN3(
        decodedPacket1_i[7]), .IN4(n528), .Q(n262) );
  AO22X1 U262 ( .IN1(decodedPacket1_o[8]), .IN2(n561), .IN3(
        decodedPacket1_i[8]), .IN4(n528), .Q(n263) );
  AO22X1 U263 ( .IN1(decodedPacket1_o[9]), .IN2(n561), .IN3(
        decodedPacket1_i[9]), .IN4(n528), .Q(n264) );
  AO22X1 U264 ( .IN1(decodedPacket1_o[10]), .IN2(n561), .IN3(
        decodedPacket1_i[10]), .IN4(n527), .Q(n265) );
  AO22X1 U265 ( .IN1(decodedPacket1_o[11]), .IN2(n561), .IN3(
        decodedPacket1_i[11]), .IN4(n527), .Q(n266) );
  AO22X1 U266 ( .IN1(decodedPacket1_o[12]), .IN2(n561), .IN3(
        decodedPacket1_i[12]), .IN4(n527), .Q(n267) );
  AO22X1 U267 ( .IN1(decodedPacket1_o[13]), .IN2(n561), .IN3(
        decodedPacket1_i[13]), .IN4(n527), .Q(n268) );
  AO22X1 U268 ( .IN1(decodedPacket1_o[14]), .IN2(n561), .IN3(
        decodedPacket1_i[14]), .IN4(n527), .Q(n269) );
  AO22X1 U269 ( .IN1(decodedPacket1_o[15]), .IN2(n561), .IN3(
        decodedPacket1_i[15]), .IN4(n527), .Q(n270) );
  AO22X1 U270 ( .IN1(decodedPacket1_o[16]), .IN2(n560), .IN3(
        decodedPacket1_i[16]), .IN4(n527), .Q(n271) );
  AO22X1 U271 ( .IN1(decodedPacket1_o[17]), .IN2(n560), .IN3(
        decodedPacket1_i[17]), .IN4(n527), .Q(n272) );
  AO22X1 U272 ( .IN1(decodedPacket1_o[18]), .IN2(n560), .IN3(
        decodedPacket1_i[18]), .IN4(n527), .Q(n273) );
  AO22X1 U273 ( .IN1(decodedPacket1_o[19]), .IN2(n560), .IN3(
        decodedPacket1_i[19]), .IN4(n527), .Q(n274) );
  AO22X1 U274 ( .IN1(decodedPacket1_o[20]), .IN2(n560), .IN3(
        decodedPacket1_i[20]), .IN4(n527), .Q(n275) );
  AO22X1 U275 ( .IN1(decodedPacket1_o[21]), .IN2(n560), .IN3(
        decodedPacket1_i[21]), .IN4(n527), .Q(n276) );
  AO22X1 U276 ( .IN1(decodedPacket1_o[22]), .IN2(n560), .IN3(
        decodedPacket1_i[22]), .IN4(n527), .Q(n277) );
  AO22X1 U277 ( .IN1(decodedPacket1_o[23]), .IN2(n560), .IN3(
        decodedPacket1_i[23]), .IN4(n527), .Q(n278) );
  AO22X1 U278 ( .IN1(decodedPacket1_o[24]), .IN2(n560), .IN3(
        decodedPacket1_i[24]), .IN4(n527), .Q(n279) );
  AO22X1 U279 ( .IN1(decodedPacket1_o[25]), .IN2(n560), .IN3(
        decodedPacket1_i[25]), .IN4(n527), .Q(n280) );
  AO22X1 U280 ( .IN1(decodedPacket1_o[26]), .IN2(n560), .IN3(
        decodedPacket1_i[26]), .IN4(n527), .Q(n281) );
  AO22X1 U281 ( .IN1(decodedPacket1_o[27]), .IN2(n560), .IN3(
        decodedPacket1_i[27]), .IN4(n527), .Q(n282) );
  AO22X1 U282 ( .IN1(decodedPacket1_o[28]), .IN2(n559), .IN3(
        decodedPacket1_i[28]), .IN4(n527), .Q(n283) );
  AO22X1 U283 ( .IN1(decodedPacket1_o[29]), .IN2(n559), .IN3(
        decodedPacket1_i[29]), .IN4(n526), .Q(n284) );
  AO22X1 U284 ( .IN1(decodedPacket1_o[30]), .IN2(n559), .IN3(
        decodedPacket1_i[30]), .IN4(n526), .Q(n285) );
  AO22X1 U285 ( .IN1(decodedPacket1_o[31]), .IN2(n559), .IN3(
        decodedPacket1_i[31]), .IN4(n526), .Q(n286) );
  AO22X1 U286 ( .IN1(decodedPacket1_o[32]), .IN2(n559), .IN3(
        decodedPacket1_i[32]), .IN4(n526), .Q(n287) );
  AO22X1 U287 ( .IN1(decodedPacket1_o[33]), .IN2(n559), .IN3(
        decodedPacket1_i[33]), .IN4(n526), .Q(n288) );
  AO22X1 U288 ( .IN1(decodedPacket1_o[34]), .IN2(n559), .IN3(
        decodedPacket1_i[34]), .IN4(n526), .Q(n289) );
  AO22X1 U289 ( .IN1(decodedPacket1_o[35]), .IN2(n559), .IN3(
        decodedPacket1_i[35]), .IN4(n526), .Q(n290) );
  AO22X1 U290 ( .IN1(decodedPacket1_o[36]), .IN2(n559), .IN3(
        decodedPacket1_i[36]), .IN4(n526), .Q(n291) );
  AO22X1 U291 ( .IN1(decodedPacket1_o[37]), .IN2(n559), .IN3(
        decodedPacket1_i[37]), .IN4(n526), .Q(n292) );
  AO22X1 U292 ( .IN1(decodedPacket1_o[38]), .IN2(n559), .IN3(
        decodedPacket1_i[38]), .IN4(n526), .Q(n293) );
  AO22X1 U293 ( .IN1(decodedPacket1_o[39]), .IN2(n559), .IN3(
        decodedPacket1_i[39]), .IN4(n526), .Q(n294) );
  AO22X1 U294 ( .IN1(decodedPacket1_o[40]), .IN2(n558), .IN3(
        decodedPacket1_i[40]), .IN4(n526), .Q(n295) );
  AO22X1 U295 ( .IN1(decodedPacket1_o[41]), .IN2(n558), .IN3(
        decodedPacket1_i[41]), .IN4(n526), .Q(n296) );
  AO22X1 U296 ( .IN1(decodedPacket1_o[42]), .IN2(n558), .IN3(
        decodedPacket1_i[42]), .IN4(n526), .Q(n297) );
  AO22X1 U297 ( .IN1(decodedPacket1_o[43]), .IN2(n558), .IN3(
        decodedPacket1_i[43]), .IN4(n526), .Q(n298) );
  AO22X1 U298 ( .IN1(decodedPacket1_o[44]), .IN2(n558), .IN3(
        decodedPacket1_i[44]), .IN4(n526), .Q(n299) );
  AO22X1 U299 ( .IN1(decodedPacket1_o[45]), .IN2(n558), .IN3(
        decodedPacket1_i[45]), .IN4(n526), .Q(n300) );
  AO22X1 U300 ( .IN1(decodedPacket1_o[46]), .IN2(n558), .IN3(
        decodedPacket1_i[46]), .IN4(n526), .Q(n301) );
  AO22X1 U301 ( .IN1(decodedPacket1_o[47]), .IN2(n558), .IN3(
        decodedPacket1_i[47]), .IN4(n526), .Q(n302) );
  AO22X1 U302 ( .IN1(decodedPacket1_o[48]), .IN2(n558), .IN3(
        decodedPacket1_i[48]), .IN4(n525), .Q(n303) );
  AO22X1 U303 ( .IN1(decodedPacket1_o[49]), .IN2(n558), .IN3(
        decodedPacket1_i[49]), .IN4(n525), .Q(n304) );
  AO22X1 U304 ( .IN1(decodedPacket1_o[50]), .IN2(n558), .IN3(
        decodedPacket1_i[50]), .IN4(n525), .Q(n305) );
  AO22X1 U305 ( .IN1(decodedPacket1_o[51]), .IN2(n558), .IN3(
        decodedPacket1_i[51]), .IN4(n525), .Q(n306) );
  AO22X1 U306 ( .IN1(decodedPacket1_o[52]), .IN2(n557), .IN3(
        decodedPacket1_i[52]), .IN4(n525), .Q(n307) );
  AO22X1 U307 ( .IN1(decodedPacket1_o[53]), .IN2(n557), .IN3(
        decodedPacket1_i[53]), .IN4(n525), .Q(n308) );
  AO22X1 U308 ( .IN1(decodedPacket1_o[54]), .IN2(n557), .IN3(
        decodedPacket1_i[54]), .IN4(n525), .Q(n309) );
  AO22X1 U309 ( .IN1(decodedPacket1_o[55]), .IN2(n557), .IN3(
        decodedPacket1_i[55]), .IN4(n525), .Q(n310) );
  AO22X1 U310 ( .IN1(decodedPacket1_o[56]), .IN2(n557), .IN3(
        decodedPacket1_i[56]), .IN4(n525), .Q(n311) );
  AO22X1 U311 ( .IN1(decodedPacket1_o[57]), .IN2(n557), .IN3(
        decodedPacket1_i[57]), .IN4(n525), .Q(n312) );
  AO22X1 U312 ( .IN1(decodedPacket1_o[58]), .IN2(n557), .IN3(
        decodedPacket1_i[58]), .IN4(n525), .Q(n313) );
  AO22X1 U313 ( .IN1(decodedPacket1_o[59]), .IN2(n557), .IN3(
        decodedPacket1_i[59]), .IN4(n525), .Q(n314) );
  AO22X1 U314 ( .IN1(decodedPacket1_o[60]), .IN2(n557), .IN3(
        decodedPacket1_i[60]), .IN4(n525), .Q(n315) );
  AO22X1 U315 ( .IN1(decodedPacket1_o[61]), .IN2(n557), .IN3(
        decodedPacket1_i[61]), .IN4(n525), .Q(n316) );
  AO22X1 U316 ( .IN1(decodedPacket1_o[62]), .IN2(n557), .IN3(
        decodedPacket1_i[62]), .IN4(n525), .Q(n317) );
  AO22X1 U317 ( .IN1(decodedPacket1_o[63]), .IN2(n557), .IN3(
        decodedPacket1_i[63]), .IN4(n525), .Q(n318) );
  AO22X1 U318 ( .IN1(decodedPacket1_o[64]), .IN2(n556), .IN3(
        decodedPacket1_i[64]), .IN4(n525), .Q(n319) );
  AO22X1 U319 ( .IN1(decodedPacket1_o[65]), .IN2(n556), .IN3(
        decodedPacket1_i[65]), .IN4(n525), .Q(n320) );
  AO22X1 U320 ( .IN1(decodedPacket1_o[66]), .IN2(n556), .IN3(
        decodedPacket1_i[66]), .IN4(n525), .Q(n321) );
  AO22X1 U321 ( .IN1(decodedPacket1_o[67]), .IN2(n556), .IN3(
        decodedPacket1_i[67]), .IN4(n524), .Q(n322) );
  AO22X1 U322 ( .IN1(decodedPacket1_o[68]), .IN2(n556), .IN3(
        decodedPacket1_i[68]), .IN4(n524), .Q(n323) );
  AO22X1 U323 ( .IN1(decodedPacket1_o[69]), .IN2(n556), .IN3(
        decodedPacket1_i[69]), .IN4(n524), .Q(n324) );
  AO22X1 U324 ( .IN1(decodedPacket1_o[70]), .IN2(n556), .IN3(
        decodedPacket1_i[70]), .IN4(n524), .Q(n325) );
  AO22X1 U325 ( .IN1(decodedPacket1_o[71]), .IN2(n556), .IN3(
        decodedPacket1_i[71]), .IN4(n524), .Q(n326) );
  AO22X1 U326 ( .IN1(decodedPacket1_o[72]), .IN2(n556), .IN3(
        decodedPacket1_i[72]), .IN4(n524), .Q(n327) );
  AO22X1 U327 ( .IN1(decodedPacket1_o[73]), .IN2(n556), .IN3(
        decodedPacket1_i[73]), .IN4(n524), .Q(n328) );
  AO22X1 U328 ( .IN1(decodedPacket1_o[74]), .IN2(n556), .IN3(
        decodedPacket1_i[74]), .IN4(n524), .Q(n329) );
  AO22X1 U329 ( .IN1(decodedPacket1_o[75]), .IN2(n556), .IN3(
        decodedPacket1_i[75]), .IN4(n524), .Q(n330) );
  AO22X1 U330 ( .IN1(decodedPacket1_o[76]), .IN2(n555), .IN3(
        decodedPacket1_i[76]), .IN4(n524), .Q(n331) );
  AO22X1 U331 ( .IN1(decodedPacket1_o[77]), .IN2(n555), .IN3(
        decodedPacket1_i[77]), .IN4(n524), .Q(n332) );
  AO22X1 U332 ( .IN1(decodedPacket1_o[78]), .IN2(n555), .IN3(
        decodedPacket1_i[78]), .IN4(n524), .Q(n333) );
  AO22X1 U333 ( .IN1(decodedPacket1_o[79]), .IN2(n555), .IN3(
        decodedPacket1_i[79]), .IN4(n524), .Q(n334) );
  AO22X1 U334 ( .IN1(decodedPacket1_o[80]), .IN2(n555), .IN3(
        decodedPacket1_i[80]), .IN4(n524), .Q(n335) );
  AO22X1 U335 ( .IN1(decodedPacket1_o[81]), .IN2(n555), .IN3(
        decodedPacket1_i[81]), .IN4(n524), .Q(n336) );
  AO22X1 U336 ( .IN1(decodedPacket1_o[82]), .IN2(n555), .IN3(
        decodedPacket1_i[82]), .IN4(n524), .Q(n337) );
  AO22X1 U337 ( .IN1(decodedPacket1_o[83]), .IN2(n555), .IN3(
        decodedPacket1_i[83]), .IN4(n524), .Q(n338) );
  AO22X1 U338 ( .IN1(decodedPacket1_o[84]), .IN2(n555), .IN3(
        decodedPacket1_i[84]), .IN4(n524), .Q(n339) );
  AO22X1 U339 ( .IN1(decodedPacket1_o[85]), .IN2(n555), .IN3(
        decodedPacket1_i[85]), .IN4(n524), .Q(n340) );
  AO22X1 U340 ( .IN1(decodedPacket1_o[86]), .IN2(n555), .IN3(
        decodedPacket1_i[86]), .IN4(n523), .Q(n341) );
  AO22X1 U341 ( .IN1(decodedPacket1_o[87]), .IN2(n555), .IN3(
        decodedPacket1_i[87]), .IN4(n523), .Q(n342) );
  AO22X1 U342 ( .IN1(decodedPacket1_o[88]), .IN2(n554), .IN3(
        decodedPacket1_i[88]), .IN4(n523), .Q(n343) );
  AO22X1 U343 ( .IN1(decodedPacket1_o[89]), .IN2(n554), .IN3(
        decodedPacket1_i[89]), .IN4(n523), .Q(n344) );
  AO22X1 U344 ( .IN1(decodedPacket1_o[90]), .IN2(n554), .IN3(
        decodedPacket1_i[90]), .IN4(n523), .Q(n345) );
  AO22X1 U345 ( .IN1(decodedPacket1_o[91]), .IN2(n554), .IN3(
        decodedPacket1_i[91]), .IN4(n523), .Q(n346) );
  AO22X1 U346 ( .IN1(decodedPacket1_o[92]), .IN2(n554), .IN3(
        decodedPacket1_i[92]), .IN4(n523), .Q(n347) );
  AO22X1 U347 ( .IN1(decodedPacket1_o[93]), .IN2(n554), .IN3(
        decodedPacket1_i[93]), .IN4(n523), .Q(n348) );
  AO22X1 U348 ( .IN1(decodedPacket1_o[94]), .IN2(n554), .IN3(
        decodedPacket1_i[94]), .IN4(n523), .Q(n349) );
  AO22X1 U349 ( .IN1(decodedPacket1_o[95]), .IN2(n554), .IN3(
        decodedPacket1_i[95]), .IN4(n523), .Q(n350) );
  AO22X1 U350 ( .IN1(decodedPacket1_o[96]), .IN2(n554), .IN3(
        decodedPacket1_i[96]), .IN4(n523), .Q(n351) );
  AO22X1 U351 ( .IN1(decodedPacket1_o[97]), .IN2(n554), .IN3(
        decodedPacket1_i[97]), .IN4(n523), .Q(n352) );
  AO22X1 U352 ( .IN1(decodedPacket1_o[98]), .IN2(n554), .IN3(
        decodedPacket1_i[98]), .IN4(n523), .Q(n353) );
  AO22X1 U353 ( .IN1(decodedPacket1_o[99]), .IN2(n554), .IN3(
        decodedPacket1_i[99]), .IN4(n523), .Q(n354) );
  AO22X1 U354 ( .IN1(decodedPacket1_o[100]), .IN2(n553), .IN3(
        decodedPacket1_i[100]), .IN4(n523), .Q(n355) );
  AO22X1 U355 ( .IN1(decodedPacket1_o[101]), .IN2(n553), .IN3(
        decodedPacket1_i[101]), .IN4(n523), .Q(n356) );
  AO22X1 U356 ( .IN1(decodedPacket1_o[102]), .IN2(n553), .IN3(
        decodedPacket1_i[102]), .IN4(n523), .Q(n357) );
  AO22X1 U357 ( .IN1(decodedPacket1_o[103]), .IN2(n553), .IN3(
        decodedPacket1_i[103]), .IN4(n523), .Q(n358) );
  AO22X1 U358 ( .IN1(decodedPacket1_o[104]), .IN2(n553), .IN3(
        decodedPacket1_i[104]), .IN4(n523), .Q(n359) );
  AO22X1 U359 ( .IN1(decodedPacket1_o[105]), .IN2(n553), .IN3(
        decodedPacket1_i[105]), .IN4(n522), .Q(n360) );
  AO22X1 U360 ( .IN1(decodedPacket1_o[106]), .IN2(n553), .IN3(
        decodedPacket1_i[106]), .IN4(n522), .Q(n361) );
  AO22X1 U361 ( .IN1(decodedPacket1_o[107]), .IN2(n553), .IN3(
        decodedPacket1_i[107]), .IN4(n522), .Q(n362) );
  AO22X1 U362 ( .IN1(decodedPacket1_o[108]), .IN2(n553), .IN3(
        decodedPacket1_i[108]), .IN4(n522), .Q(n363) );
  AO22X1 U363 ( .IN1(decodedPacket1_o[109]), .IN2(n553), .IN3(
        decodedPacket1_i[109]), .IN4(n522), .Q(n364) );
  AO22X1 U364 ( .IN1(decodedPacket1_o[110]), .IN2(n553), .IN3(
        decodedPacket1_i[110]), .IN4(n522), .Q(n365) );
  AO22X1 U365 ( .IN1(decodedPacket1_o[111]), .IN2(n553), .IN3(
        decodedPacket1_i[111]), .IN4(n522), .Q(n366) );
  AO22X1 U366 ( .IN1(decodedPacket1_o[112]), .IN2(n552), .IN3(
        decodedPacket1_i[112]), .IN4(n522), .Q(n367) );
  AO22X1 U367 ( .IN1(decodedPacket1_o[113]), .IN2(n552), .IN3(
        decodedPacket1_i[113]), .IN4(n522), .Q(n368) );
  AO22X1 U368 ( .IN1(decodedPacket1_o[114]), .IN2(n552), .IN3(
        decodedPacket1_i[114]), .IN4(n522), .Q(n369) );
  AO22X1 U369 ( .IN1(decodedPacket1_o[115]), .IN2(n552), .IN3(
        decodedPacket1_i[115]), .IN4(n522), .Q(n370) );
  AO22X1 U370 ( .IN1(decodedPacket1_o[116]), .IN2(n552), .IN3(
        decodedPacket1_i[116]), .IN4(n522), .Q(n371) );
  AO22X1 U371 ( .IN1(decodedPacket1_o[117]), .IN2(n552), .IN3(
        decodedPacket1_i[117]), .IN4(n522), .Q(n372) );
  AO22X1 U372 ( .IN1(decodedPacket1_o[118]), .IN2(n552), .IN3(
        decodedPacket1_i[118]), .IN4(n522), .Q(n373) );
  AO22X1 U373 ( .IN1(decodedPacket1_o[119]), .IN2(n552), .IN3(
        decodedPacket1_i[119]), .IN4(n522), .Q(n374) );
  AO22X1 U374 ( .IN1(decodedPacket1_o[120]), .IN2(n552), .IN3(
        decodedPacket1_i[120]), .IN4(n522), .Q(n375) );
  AO22X1 U375 ( .IN1(decodedPacket1_o[121]), .IN2(n552), .IN3(
        decodedPacket1_i[121]), .IN4(n522), .Q(n376) );
  AO22X1 U376 ( .IN1(decodedPacket1_o[122]), .IN2(n552), .IN3(
        decodedPacket1_i[122]), .IN4(n522), .Q(n377) );
  AO22X1 U377 ( .IN1(decodedPacket1_o[123]), .IN2(n552), .IN3(
        decodedPacket1_i[123]), .IN4(n522), .Q(n378) );
  AO22X1 U378 ( .IN1(decodedPacket1_o[124]), .IN2(n551), .IN3(
        decodedPacket1_i[124]), .IN4(n521), .Q(n379) );
  AO22X1 U379 ( .IN1(decodedPacket1_o[125]), .IN2(n551), .IN3(
        decodedPacket1_i[125]), .IN4(n521), .Q(n380) );
  AO22X1 U380 ( .IN1(decodedPacket0_o[0]), .IN2(n551), .IN3(
        decodedPacket0_i[0]), .IN4(n521), .Q(n381) );
  AO22X1 U381 ( .IN1(decodedPacket0_o[1]), .IN2(n551), .IN3(
        decodedPacket0_i[1]), .IN4(n521), .Q(n382) );
  AO22X1 U382 ( .IN1(decodedPacket0_o[2]), .IN2(n551), .IN3(
        decodedPacket0_i[2]), .IN4(n521), .Q(n383) );
  AO22X1 U383 ( .IN1(decodedPacket0_o[3]), .IN2(n551), .IN3(
        decodedPacket0_i[3]), .IN4(n521), .Q(n384) );
  AO22X1 U384 ( .IN1(decodedPacket0_o[4]), .IN2(n551), .IN3(
        decodedPacket0_i[4]), .IN4(n521), .Q(n385) );
  AO22X1 U385 ( .IN1(decodedPacket0_o[5]), .IN2(n551), .IN3(
        decodedPacket0_i[5]), .IN4(n521), .Q(n386) );
  AO22X1 U386 ( .IN1(decodedPacket0_o[6]), .IN2(n551), .IN3(
        decodedPacket0_i[6]), .IN4(n521), .Q(n387) );
  AO22X1 U387 ( .IN1(decodedPacket0_o[7]), .IN2(n551), .IN3(
        decodedPacket0_i[7]), .IN4(n521), .Q(n388) );
  AO22X1 U388 ( .IN1(decodedPacket0_o[8]), .IN2(n551), .IN3(
        decodedPacket0_i[8]), .IN4(n521), .Q(n389) );
  AO22X1 U389 ( .IN1(decodedPacket0_o[9]), .IN2(n551), .IN3(
        decodedPacket0_i[9]), .IN4(n521), .Q(n390) );
  AO22X1 U390 ( .IN1(decodedPacket0_o[10]), .IN2(n550), .IN3(
        decodedPacket0_i[10]), .IN4(n521), .Q(n391) );
  AO22X1 U391 ( .IN1(decodedPacket0_o[11]), .IN2(n550), .IN3(
        decodedPacket0_i[11]), .IN4(n521), .Q(n392) );
  AO22X1 U392 ( .IN1(decodedPacket0_o[12]), .IN2(n550), .IN3(
        decodedPacket0_i[12]), .IN4(n521), .Q(n393) );
  AO22X1 U393 ( .IN1(decodedPacket0_o[13]), .IN2(n550), .IN3(
        decodedPacket0_i[13]), .IN4(n521), .Q(n394) );
  AO22X1 U394 ( .IN1(decodedPacket0_o[14]), .IN2(n550), .IN3(
        decodedPacket0_i[14]), .IN4(n521), .Q(n395) );
  AO22X1 U395 ( .IN1(decodedPacket0_o[15]), .IN2(n550), .IN3(
        decodedPacket0_i[15]), .IN4(n521), .Q(n396) );
  AO22X1 U396 ( .IN1(decodedPacket0_o[16]), .IN2(n550), .IN3(
        decodedPacket0_i[16]), .IN4(n521), .Q(n397) );
  AO22X1 U397 ( .IN1(decodedPacket0_o[17]), .IN2(n550), .IN3(
        decodedPacket0_i[17]), .IN4(n520), .Q(n398) );
  AO22X1 U398 ( .IN1(decodedPacket0_o[18]), .IN2(n550), .IN3(
        decodedPacket0_i[18]), .IN4(n520), .Q(n399) );
  AO22X1 U399 ( .IN1(decodedPacket0_o[19]), .IN2(n550), .IN3(
        decodedPacket0_i[19]), .IN4(n520), .Q(n400) );
  AO22X1 U400 ( .IN1(decodedPacket0_o[20]), .IN2(n550), .IN3(
        decodedPacket0_i[20]), .IN4(n520), .Q(n401) );
  AO22X1 U401 ( .IN1(decodedPacket0_o[21]), .IN2(n550), .IN3(
        decodedPacket0_i[21]), .IN4(n520), .Q(n402) );
  AO22X1 U402 ( .IN1(decodedPacket0_o[22]), .IN2(n549), .IN3(
        decodedPacket0_i[22]), .IN4(n520), .Q(n403) );
  AO22X1 U403 ( .IN1(decodedPacket0_o[23]), .IN2(n549), .IN3(
        decodedPacket0_i[23]), .IN4(n520), .Q(n404) );
  AO22X1 U404 ( .IN1(decodedPacket0_o[24]), .IN2(n549), .IN3(
        decodedPacket0_i[24]), .IN4(n520), .Q(n405) );
  AO22X1 U405 ( .IN1(decodedPacket0_o[25]), .IN2(n549), .IN3(
        decodedPacket0_i[25]), .IN4(n520), .Q(n406) );
  AO22X1 U406 ( .IN1(decodedPacket0_o[26]), .IN2(n549), .IN3(
        decodedPacket0_i[26]), .IN4(n520), .Q(n407) );
  AO22X1 U407 ( .IN1(decodedPacket0_o[27]), .IN2(n549), .IN3(
        decodedPacket0_i[27]), .IN4(n520), .Q(n408) );
  AO22X1 U408 ( .IN1(decodedPacket0_o[28]), .IN2(n549), .IN3(
        decodedPacket0_i[28]), .IN4(n520), .Q(n409) );
  AO22X1 U409 ( .IN1(decodedPacket0_o[29]), .IN2(n549), .IN3(
        decodedPacket0_i[29]), .IN4(n520), .Q(n410) );
  AO22X1 U410 ( .IN1(decodedPacket0_o[30]), .IN2(n549), .IN3(
        decodedPacket0_i[30]), .IN4(n520), .Q(n411) );
  AO22X1 U411 ( .IN1(decodedPacket0_o[31]), .IN2(n549), .IN3(
        decodedPacket0_i[31]), .IN4(n520), .Q(n412) );
  AO22X1 U412 ( .IN1(decodedPacket0_o[32]), .IN2(n549), .IN3(
        decodedPacket0_i[32]), .IN4(n520), .Q(n413) );
  AO22X1 U413 ( .IN1(decodedPacket0_o[33]), .IN2(n549), .IN3(
        decodedPacket0_i[33]), .IN4(n520), .Q(n414) );
  AO22X1 U414 ( .IN1(decodedPacket0_o[34]), .IN2(n548), .IN3(
        decodedPacket0_i[34]), .IN4(n520), .Q(n415) );
  AO22X1 U415 ( .IN1(decodedPacket0_o[35]), .IN2(n548), .IN3(
        decodedPacket0_i[35]), .IN4(n520), .Q(n416) );
  AO22X1 U416 ( .IN1(decodedPacket0_o[36]), .IN2(n548), .IN3(
        decodedPacket0_i[36]), .IN4(n519), .Q(n417) );
  AO22X1 U417 ( .IN1(decodedPacket0_o[37]), .IN2(n548), .IN3(
        decodedPacket0_i[37]), .IN4(n519), .Q(n418) );
  AO22X1 U418 ( .IN1(decodedPacket0_o[38]), .IN2(n548), .IN3(
        decodedPacket0_i[38]), .IN4(n519), .Q(n419) );
  AO22X1 U419 ( .IN1(decodedPacket0_o[39]), .IN2(n548), .IN3(
        decodedPacket0_i[39]), .IN4(n519), .Q(n420) );
  AO22X1 U420 ( .IN1(decodedPacket0_o[40]), .IN2(n548), .IN3(
        decodedPacket0_i[40]), .IN4(n519), .Q(n421) );
  AO22X1 U421 ( .IN1(decodedPacket0_o[41]), .IN2(n548), .IN3(
        decodedPacket0_i[41]), .IN4(n519), .Q(n422) );
  AO22X1 U422 ( .IN1(decodedPacket0_o[42]), .IN2(n548), .IN3(
        decodedPacket0_i[42]), .IN4(n519), .Q(n423) );
  AO22X1 U423 ( .IN1(decodedPacket0_o[43]), .IN2(n548), .IN3(
        decodedPacket0_i[43]), .IN4(n519), .Q(n424) );
  AO22X1 U424 ( .IN1(decodedPacket0_o[44]), .IN2(n548), .IN3(
        decodedPacket0_i[44]), .IN4(n519), .Q(n425) );
  AO22X1 U425 ( .IN1(decodedPacket0_o[45]), .IN2(n548), .IN3(
        decodedPacket0_i[45]), .IN4(n519), .Q(n426) );
  AO22X1 U426 ( .IN1(decodedPacket0_o[46]), .IN2(n547), .IN3(
        decodedPacket0_i[46]), .IN4(n519), .Q(n427) );
  AO22X1 U427 ( .IN1(decodedPacket0_o[47]), .IN2(n547), .IN3(
        decodedPacket0_i[47]), .IN4(n519), .Q(n428) );
  AO22X1 U428 ( .IN1(decodedPacket0_o[48]), .IN2(n547), .IN3(
        decodedPacket0_i[48]), .IN4(n519), .Q(n429) );
  AO22X1 U429 ( .IN1(decodedPacket0_o[49]), .IN2(n547), .IN3(
        decodedPacket0_i[49]), .IN4(n519), .Q(n430) );
  AO22X1 U430 ( .IN1(decodedPacket0_o[50]), .IN2(n547), .IN3(
        decodedPacket0_i[50]), .IN4(n519), .Q(n431) );
  AO22X1 U431 ( .IN1(decodedPacket0_o[51]), .IN2(n547), .IN3(
        decodedPacket0_i[51]), .IN4(n519), .Q(n432) );
  AO22X1 U432 ( .IN1(decodedPacket0_o[52]), .IN2(n547), .IN3(
        decodedPacket0_i[52]), .IN4(n519), .Q(n433) );
  AO22X1 U433 ( .IN1(decodedPacket0_o[53]), .IN2(n547), .IN3(
        decodedPacket0_i[53]), .IN4(n519), .Q(n434) );
  AO22X1 U434 ( .IN1(decodedPacket0_o[54]), .IN2(n547), .IN3(
        decodedPacket0_i[54]), .IN4(n519), .Q(n435) );
  AO22X1 U435 ( .IN1(decodedPacket0_o[55]), .IN2(n547), .IN3(
        decodedPacket0_i[55]), .IN4(n518), .Q(n436) );
  AO22X1 U436 ( .IN1(decodedPacket0_o[56]), .IN2(n547), .IN3(
        decodedPacket0_i[56]), .IN4(n518), .Q(n437) );
  AO22X1 U437 ( .IN1(decodedPacket0_o[57]), .IN2(n547), .IN3(
        decodedPacket0_i[57]), .IN4(n518), .Q(n438) );
  AO22X1 U438 ( .IN1(decodedPacket0_o[58]), .IN2(n546), .IN3(
        decodedPacket0_i[58]), .IN4(n518), .Q(n439) );
  AO22X1 U439 ( .IN1(decodedPacket0_o[59]), .IN2(n546), .IN3(
        decodedPacket0_i[59]), .IN4(n518), .Q(n440) );
  AO22X1 U440 ( .IN1(decodedPacket0_o[60]), .IN2(n546), .IN3(
        decodedPacket0_i[60]), .IN4(n518), .Q(n441) );
  AO22X1 U441 ( .IN1(decodedPacket0_o[61]), .IN2(n546), .IN3(
        decodedPacket0_i[61]), .IN4(n518), .Q(n442) );
  AO22X1 U442 ( .IN1(decodedPacket0_o[62]), .IN2(n546), .IN3(
        decodedPacket0_i[62]), .IN4(n518), .Q(n443) );
  AO22X1 U443 ( .IN1(decodedPacket0_o[63]), .IN2(n546), .IN3(
        decodedPacket0_i[63]), .IN4(n518), .Q(n444) );
  AO22X1 U444 ( .IN1(decodedPacket0_o[64]), .IN2(n546), .IN3(
        decodedPacket0_i[64]), .IN4(n518), .Q(n445) );
  AO22X1 U445 ( .IN1(decodedPacket0_o[65]), .IN2(n546), .IN3(
        decodedPacket0_i[65]), .IN4(n518), .Q(n446) );
  AO22X1 U446 ( .IN1(decodedPacket0_o[66]), .IN2(n546), .IN3(
        decodedPacket0_i[66]), .IN4(n518), .Q(n447) );
  AO22X1 U447 ( .IN1(decodedPacket0_o[67]), .IN2(n546), .IN3(
        decodedPacket0_i[67]), .IN4(n518), .Q(n448) );
  AO22X1 U448 ( .IN1(decodedPacket0_o[68]), .IN2(n546), .IN3(
        decodedPacket0_i[68]), .IN4(n518), .Q(n449) );
  AO22X1 U449 ( .IN1(decodedPacket0_o[69]), .IN2(n546), .IN3(
        decodedPacket0_i[69]), .IN4(n518), .Q(n450) );
  AO22X1 U450 ( .IN1(decodedPacket0_o[70]), .IN2(n545), .IN3(
        decodedPacket0_i[70]), .IN4(n518), .Q(n451) );
  AO22X1 U451 ( .IN1(decodedPacket0_o[71]), .IN2(n545), .IN3(
        decodedPacket0_i[71]), .IN4(n518), .Q(n452) );
  AO22X1 U452 ( .IN1(decodedPacket0_o[72]), .IN2(n545), .IN3(
        decodedPacket0_i[72]), .IN4(n518), .Q(n453) );
  AO22X1 U453 ( .IN1(decodedPacket0_o[73]), .IN2(n545), .IN3(
        decodedPacket0_i[73]), .IN4(n518), .Q(n454) );
  AO22X1 U454 ( .IN1(decodedPacket0_o[74]), .IN2(n545), .IN3(
        decodedPacket0_i[74]), .IN4(n512), .Q(n455) );
  AO22X1 U455 ( .IN1(decodedPacket0_o[75]), .IN2(n545), .IN3(
        decodedPacket0_i[75]), .IN4(n512), .Q(n456) );
  AO22X1 U456 ( .IN1(decodedPacket0_o[76]), .IN2(n545), .IN3(
        decodedPacket0_i[76]), .IN4(n515), .Q(n457) );
  AO22X1 U457 ( .IN1(decodedPacket0_o[77]), .IN2(n545), .IN3(
        decodedPacket0_i[77]), .IN4(n514), .Q(n458) );
  AO22X1 U458 ( .IN1(decodedPacket0_o[78]), .IN2(n545), .IN3(
        decodedPacket0_i[78]), .IN4(n511), .Q(n459) );
  AO22X1 U459 ( .IN1(decodedPacket0_o[79]), .IN2(n545), .IN3(
        decodedPacket0_i[79]), .IN4(n513), .Q(n460) );
  AO22X1 U460 ( .IN1(decodedPacket0_o[80]), .IN2(n545), .IN3(
        decodedPacket0_i[80]), .IN4(n529), .Q(n461) );
  AO22X1 U461 ( .IN1(decodedPacket0_o[81]), .IN2(n545), .IN3(
        decodedPacket0_i[81]), .IN4(n516), .Q(n462) );
  AO22X1 U462 ( .IN1(decodedPacket0_o[82]), .IN2(n544), .IN3(
        decodedPacket0_i[82]), .IN4(n524), .Q(n463) );
  AO22X1 U463 ( .IN1(decodedPacket0_o[83]), .IN2(n544), .IN3(
        decodedPacket0_i[83]), .IN4(n512), .Q(n464) );
  AO22X1 U464 ( .IN1(decodedPacket0_o[84]), .IN2(n544), .IN3(
        decodedPacket0_i[84]), .IN4(n515), .Q(n465) );
  AO22X1 U465 ( .IN1(decodedPacket0_o[85]), .IN2(n544), .IN3(
        decodedPacket0_i[85]), .IN4(n514), .Q(n466) );
  AO22X1 U466 ( .IN1(decodedPacket0_o[86]), .IN2(n544), .IN3(
        decodedPacket0_i[86]), .IN4(n511), .Q(n467) );
  AO22X1 U467 ( .IN1(decodedPacket0_o[87]), .IN2(n544), .IN3(
        decodedPacket0_i[87]), .IN4(n513), .Q(n468) );
  AO22X1 U468 ( .IN1(decodedPacket0_o[88]), .IN2(n544), .IN3(
        decodedPacket0_i[88]), .IN4(n516), .Q(n469) );
  AO22X1 U469 ( .IN1(decodedPacket0_o[89]), .IN2(n544), .IN3(
        decodedPacket0_i[89]), .IN4(n516), .Q(n470) );
  AO22X1 U470 ( .IN1(decodedPacket0_o[90]), .IN2(n544), .IN3(
        decodedPacket0_i[90]), .IN4(n525), .Q(n471) );
  AO22X1 U471 ( .IN1(decodedPacket0_o[91]), .IN2(n544), .IN3(
        decodedPacket0_i[91]), .IN4(n512), .Q(n472) );
  AO22X1 U472 ( .IN1(decodedPacket0_o[92]), .IN2(n544), .IN3(
        decodedPacket0_i[92]), .IN4(n515), .Q(n473) );
  AO22X1 U473 ( .IN1(decodedPacket0_o[93]), .IN2(n544), .IN3(
        decodedPacket0_i[93]), .IN4(n517), .Q(n474) );
  AO22X1 U474 ( .IN1(decodedPacket0_o[94]), .IN2(n543), .IN3(
        decodedPacket0_i[94]), .IN4(n517), .Q(n475) );
  AO22X1 U475 ( .IN1(decodedPacket0_o[95]), .IN2(n543), .IN3(
        decodedPacket0_i[95]), .IN4(n517), .Q(n476) );
  AO22X1 U476 ( .IN1(decodedPacket0_o[96]), .IN2(n543), .IN3(
        decodedPacket0_i[96]), .IN4(n517), .Q(n477) );
  AO22X1 U477 ( .IN1(decodedPacket0_o[97]), .IN2(n543), .IN3(
        decodedPacket0_i[97]), .IN4(n517), .Q(n478) );
  AO22X1 U478 ( .IN1(decodedPacket0_o[98]), .IN2(n543), .IN3(
        decodedPacket0_i[98]), .IN4(n517), .Q(n479) );
  AO22X1 U479 ( .IN1(decodedPacket0_o[99]), .IN2(n543), .IN3(
        decodedPacket0_i[99]), .IN4(n517), .Q(n480) );
  AO22X1 U480 ( .IN1(decodedPacket0_o[100]), .IN2(n543), .IN3(
        decodedPacket0_i[100]), .IN4(n517), .Q(n481) );
  AO22X1 U481 ( .IN1(decodedPacket0_o[101]), .IN2(n543), .IN3(
        decodedPacket0_i[101]), .IN4(n517), .Q(n482) );
  AO22X1 U482 ( .IN1(decodedPacket0_o[102]), .IN2(n543), .IN3(
        decodedPacket0_i[102]), .IN4(n517), .Q(n483) );
  AO22X1 U483 ( .IN1(decodedPacket0_o[103]), .IN2(n543), .IN3(
        decodedPacket0_i[103]), .IN4(n517), .Q(n484) );
  AO22X1 U484 ( .IN1(decodedPacket0_o[104]), .IN2(n543), .IN3(
        decodedPacket0_i[104]), .IN4(n517), .Q(n485) );
  AO22X1 U485 ( .IN1(decodedPacket0_o[105]), .IN2(n543), .IN3(
        decodedPacket0_i[105]), .IN4(n517), .Q(n486) );
  AO22X1 U486 ( .IN1(decodedPacket0_o[106]), .IN2(n542), .IN3(
        decodedPacket0_i[106]), .IN4(n517), .Q(n487) );
  AO22X1 U487 ( .IN1(decodedPacket0_o[107]), .IN2(n542), .IN3(
        decodedPacket0_i[107]), .IN4(n517), .Q(n488) );
  AO22X1 U488 ( .IN1(decodedPacket0_o[108]), .IN2(n542), .IN3(
        decodedPacket0_i[108]), .IN4(n517), .Q(n489) );
  AO22X1 U489 ( .IN1(decodedPacket0_o[109]), .IN2(n542), .IN3(
        decodedPacket0_i[109]), .IN4(n517), .Q(n490) );
  AO22X1 U490 ( .IN1(decodedPacket0_o[110]), .IN2(n542), .IN3(
        decodedPacket0_i[110]), .IN4(n517), .Q(n491) );
  AO22X1 U491 ( .IN1(decodedPacket0_o[111]), .IN2(n542), .IN3(
        decodedPacket0_i[111]), .IN4(n517), .Q(n492) );
  AO22X1 U492 ( .IN1(decodedPacket0_o[112]), .IN2(n542), .IN3(
        decodedPacket0_i[112]), .IN4(n540), .Q(n493) );
  AO22X1 U493 ( .IN1(decodedPacket0_o[113]), .IN2(n542), .IN3(
        decodedPacket0_i[113]), .IN4(n540), .Q(n494) );
  AO22X1 U494 ( .IN1(decodedPacket0_o[114]), .IN2(n542), .IN3(
        decodedPacket0_i[114]), .IN4(n540), .Q(n495) );
  AO22X1 U495 ( .IN1(decodedPacket0_o[115]), .IN2(n542), .IN3(
        decodedPacket0_i[115]), .IN4(n511), .Q(n496) );
  AO22X1 U496 ( .IN1(decodedPacket0_o[116]), .IN2(n542), .IN3(
        decodedPacket0_i[116]), .IN4(n540), .Q(n497) );
  AO22X1 U497 ( .IN1(decodedPacket0_o[117]), .IN2(n542), .IN3(
        decodedPacket0_i[117]), .IN4(n511), .Q(n498) );
  AO22X1 U498 ( .IN1(decodedPacket0_o[118]), .IN2(n541), .IN3(
        decodedPacket0_i[118]), .IN4(n516), .Q(n499) );
  AO22X1 U499 ( .IN1(decodedPacket0_o[119]), .IN2(n541), .IN3(
        decodedPacket0_i[119]), .IN4(n515), .Q(n500) );
  AO22X1 U500 ( .IN1(decodedPacket0_o[120]), .IN2(n541), .IN3(
        decodedPacket0_i[120]), .IN4(n514), .Q(n501) );
  AO22X1 U501 ( .IN1(decodedPacket0_o[121]), .IN2(n541), .IN3(
        decodedPacket0_i[121]), .IN4(n526), .Q(n502) );
  AO22X1 U502 ( .IN1(decodedPacket0_o[122]), .IN2(n541), .IN3(
        decodedPacket0_i[122]), .IN4(n512), .Q(n503) );
  AO22X1 U503 ( .IN1(decodedPacket0_o[123]), .IN2(n541), .IN3(
        decodedPacket0_i[123]), .IN4(n511), .Q(n504) );
  AO22X1 U504 ( .IN1(decodedPacket0_o[124]), .IN2(n541), .IN3(
        decodedPacket0_i[124]), .IN4(n511), .Q(n505) );
  AO22X1 U505 ( .IN1(decodedPacket0_o[125]), .IN2(n541), .IN3(
        decodedPacket0_i[125]), .IN4(n513), .Q(n506) );
  AO22X1 U506 ( .IN1(instBufferReady_o), .IN2(n541), .IN3(instBufferReady_i), 
        .IN4(n513), .Q(n507) );
  AO22X1 U507 ( .IN1(branchCount_o[0]), .IN2(n541), .IN3(branchCount_i[0]), 
        .IN4(n516), .Q(n508) );
  AO22X1 U508 ( .IN1(branchCount_o[1]), .IN2(n541), .IN3(branchCount_i[1]), 
        .IN4(n515), .Q(n509) );
  AO22X1 U509 ( .IN1(branchCount_o[2]), .IN2(n541), .IN3(branchCount_i[2]), 
        .IN4(n514), .Q(n510) );
  NOR3X0 U510 ( .IN1(flush_i), .IN2(reset), .IN3(n2), .QN(n1) );
  NOR3X0 U511 ( .IN1(stall_i), .IN2(reset), .IN3(flush_i), .QN(n2) );
  NBUFFX2 U512 ( .INP(n578), .Z(n572) );
  NBUFFX2 U513 ( .INP(n578), .Z(n571) );
  NBUFFX2 U514 ( .INP(n580), .Z(n562) );
  NBUFFX2 U515 ( .INP(n578), .Z(n561) );
  NBUFFX2 U516 ( .INP(n580), .Z(n560) );
  NBUFFX2 U517 ( .INP(n579), .Z(n550) );
  NBUFFX2 U518 ( .INP(n579), .Z(n549) );
  NBUFFX2 U519 ( .INP(n579), .Z(n548) );
  NBUFFX2 U520 ( .INP(n578), .Z(n577) );
  NBUFFX2 U521 ( .INP(n1), .Z(n564) );
  NBUFFX2 U522 ( .INP(n1), .Z(n563) );
  NBUFFX2 U523 ( .INP(n579), .Z(n553) );
  NBUFFX2 U524 ( .INP(n579), .Z(n552) );
  NBUFFX2 U525 ( .INP(n579), .Z(n551) );
  NBUFFX2 U526 ( .INP(n1), .Z(n580) );
  NBUFFX2 U527 ( .INP(n2), .Z(n516) );
  NBUFFX2 U528 ( .INP(n2), .Z(n515) );
  NBUFFX2 U529 ( .INP(n2), .Z(n514) );
  NBUFFX2 U530 ( .INP(n2), .Z(n513) );
  NBUFFX2 U531 ( .INP(n2), .Z(n512) );
  NBUFFX2 U532 ( .INP(n2), .Z(n511) );
  NBUFFX2 U533 ( .INP(n514), .Z(n517) );
  NBUFFX2 U534 ( .INP(n511), .Z(n518) );
  NBUFFX2 U535 ( .INP(n511), .Z(n519) );
  NBUFFX2 U536 ( .INP(n511), .Z(n520) );
  NBUFFX2 U537 ( .INP(n512), .Z(n521) );
  NBUFFX2 U538 ( .INP(n512), .Z(n522) );
  NBUFFX2 U539 ( .INP(n512), .Z(n523) );
  NBUFFX2 U540 ( .INP(n513), .Z(n524) );
  NBUFFX2 U541 ( .INP(n513), .Z(n525) );
  NBUFFX2 U542 ( .INP(n513), .Z(n526) );
  NBUFFX2 U543 ( .INP(n512), .Z(n527) );
  NBUFFX2 U544 ( .INP(n513), .Z(n528) );
  NBUFFX2 U545 ( .INP(n515), .Z(n529) );
  NBUFFX2 U546 ( .INP(n514), .Z(n530) );
  NBUFFX2 U547 ( .INP(n514), .Z(n531) );
  NBUFFX2 U548 ( .INP(n514), .Z(n532) );
  NBUFFX2 U549 ( .INP(n515), .Z(n533) );
  NBUFFX2 U550 ( .INP(n515), .Z(n534) );
  NBUFFX2 U551 ( .INP(n515), .Z(n535) );
  NBUFFX2 U552 ( .INP(n516), .Z(n536) );
  NBUFFX2 U553 ( .INP(n516), .Z(n537) );
  NBUFFX2 U554 ( .INP(n514), .Z(n538) );
  NBUFFX2 U555 ( .INP(n512), .Z(n539) );
  NBUFFX2 U556 ( .INP(n515), .Z(n540) );
  NBUFFX2 U557 ( .INP(n580), .Z(n541) );
  NBUFFX2 U558 ( .INP(n580), .Z(n542) );
  NBUFFX2 U559 ( .INP(n580), .Z(n543) );
  NBUFFX2 U560 ( .INP(n580), .Z(n544) );
  NBUFFX2 U561 ( .INP(n580), .Z(n545) );
  NBUFFX2 U562 ( .INP(n580), .Z(n546) );
  NBUFFX2 U563 ( .INP(n580), .Z(n547) );
  NBUFFX2 U564 ( .INP(n579), .Z(n554) );
  NBUFFX2 U565 ( .INP(n579), .Z(n555) );
  NBUFFX2 U566 ( .INP(n579), .Z(n556) );
  NBUFFX2 U567 ( .INP(n579), .Z(n557) );
  NBUFFX2 U568 ( .INP(n579), .Z(n558) );
  NBUFFX2 U569 ( .INP(n579), .Z(n559) );
  NBUFFX2 U570 ( .INP(n1), .Z(n565) );
  NBUFFX2 U571 ( .INP(n1), .Z(n566) );
  NBUFFX2 U572 ( .INP(n1), .Z(n567) );
  NBUFFX2 U573 ( .INP(n1), .Z(n568) );
  NBUFFX2 U574 ( .INP(n1), .Z(n569) );
  NBUFFX2 U575 ( .INP(n1), .Z(n570) );
  NBUFFX2 U576 ( .INP(n578), .Z(n573) );
  NBUFFX2 U577 ( .INP(n578), .Z(n574) );
  NBUFFX2 U578 ( .INP(n578), .Z(n575) );
  NBUFFX2 U579 ( .INP(n578), .Z(n576) );
  NBUFFX2 U580 ( .INP(n1), .Z(n578) );
  NBUFFX2 U581 ( .INP(n1), .Z(n579) );
endmodule

