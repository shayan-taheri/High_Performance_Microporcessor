
module Dispatch ( clk, reset, stall_i, renameReady_i, flagRecoverEX_i, 
        ctrlVerified_i, ctrlVerifiedSMTid_i, renamedPacket0_i, 
        renamedPacket1_i, renamedPacket2_i, renamedPacket3_i, loadQueueCnt_i, 
        storeQueueCnt_i, issueQueueCnt_i, activeListCnt_i, issueqPacket0_o, 
        issueqPacket1_o, issueqPacket2_o, issueqPacket3_o, alPacket0_o, 
        alPacket1_o, alPacket2_o, alPacket3_o, lsqPacket0_o, lsqPacket1_o, 
        lsqPacket2_o, lsqPacket3_o, updatedBranchMask0_o, updatedBranchMask1_o, 
        updatedBranchMask2_o, updatedBranchMask3_o, backEndReady_o, 
        stallfrontEnd_o );
  input [1:0] ctrlVerifiedSMTid_i;
  input [144:0] renamedPacket0_i;
  input [144:0] renamedPacket1_i;
  input [144:0] renamedPacket2_i;
  input [144:0] renamedPacket3_i;
  input [5:0] loadQueueCnt_i;
  input [5:0] storeQueueCnt_i;
  input [5:0] issueQueueCnt_i;
  input [7:0] activeListCnt_i;
  output [144:0] issueqPacket0_o;
  output [144:0] issueqPacket1_o;
  output [144:0] issueqPacket2_o;
  output [144:0] issueqPacket3_o;
  output [54:0] alPacket0_o;
  output [54:0] alPacket1_o;
  output [54:0] alPacket2_o;
  output [54:0] alPacket3_o;
  output [5:0] lsqPacket0_o;
  output [5:0] lsqPacket1_o;
  output [5:0] lsqPacket2_o;
  output [5:0] lsqPacket3_o;
  output [3:0] updatedBranchMask0_o;
  output [3:0] updatedBranchMask1_o;
  output [3:0] updatedBranchMask2_o;
  output [3:0] updatedBranchMask3_o;
  input clk, reset, stall_i, renameReady_i, flagRecoverEX_i, ctrlVerified_i;
  output backEndReady_o, stallfrontEnd_o;
  wire   issueqPacket0_o_138, issueqPacket0_o_131, issueqPacket0_o_130,
         issueqPacket0_o_122, issueqPacket0_o_36, issueqPacket0_o_35,
         issueqPacket0_o_34, issueqPacket0_o_33, issueqPacket0_o_32,
         issueqPacket0_o_31, issueqPacket0_o_30, issueqPacket0_o_29,
         issueqPacket0_o_28, issueqPacket0_o_27, issueqPacket0_o_26,
         issueqPacket0_o_25, issueqPacket0_o_24, issueqPacket0_o_23,
         issueqPacket0_o_22, issueqPacket0_o_21, issueqPacket0_o_20,
         issueqPacket0_o_19, issueqPacket0_o_18, issueqPacket0_o_17,
         issueqPacket0_o_16, issueqPacket0_o_15, issueqPacket0_o_14,
         issueqPacket0_o_13, issueqPacket0_o_12, issueqPacket0_o_11,
         issueqPacket0_o_10, issueqPacket0_o_9, issueqPacket0_o_8,
         issueqPacket0_o_7, issueqPacket0_o_6, issueqPacket0_o_5,
         issueqPacket0_o_4, issueqPacket0_o_3, issueqPacket0_o_2,
         issueqPacket0_o_1, issueqPacket0_o_0, issueqPacket1_o_144,
         issueqPacket1_o_143, issueqPacket1_o_142, issueqPacket1_o_141,
         issueqPacket1_o_140, issueqPacket1_o_139, issueqPacket1_o_138,
         issueqPacket1_o_137, issueqPacket1_o_136, issueqPacket2_o_144,
         issueqPacket2_o_143, issueqPacket2_o_142, issueqPacket2_o_141,
         issueqPacket2_o_140, issueqPacket2_o_139, issueqPacket2_o_138,
         issueqPacket2_o_137, issueqPacket2_o_136, issueqPacket3_o_144,
         issueqPacket3_o_143, issueqPacket3_o_142, issueqPacket3_o_141,
         issueqPacket3_o_140, issueqPacket3_o_139, issueqPacket3_o_138, N22,
         N23, N24, N25, N26, N27, N28, stall0, N29, N30, N31, N32, N33, N34,
         N35, stall1, stall2, stall3, N51, N50, N49, N48, N47, N46, N45, N44,
         N43, N42, N41, N40, N39, N38, N37, N36, n61, n62, n63, n64, n65,
         \loadCnt[2] , \loadCnt[1] , \loadCnt[0] , N5, N4, \storeCnt[2] ,
         \storeCnt[1] , \storeCnt[0] , N9, N10, \add_291/carry[7] ,
         \add_291/carry[6] , \add_291/carry[5] , \add_291/carry[4] ,
         \add_290/carry[5] , \add_290/carry[4] , \add_288/carry[5] ,
         \add_288/carry[4] , \add_288/carry[3] , \add_288/carry[2] ,
         \add_288/carry[1] , \add_289/carry[5] , \add_289/carry[4] ,
         \add_289/carry[3] , \add_289/carry[2] , \add_289/carry[1] , n66, n69,
         n72, n75, n78, n81, n84, n87, n90, n93, n96, n99, n102, n105, n108,
         n111, n114, n118, n122, n125, n128, n131, n134, n137, n140, n143,
         n146, n149, n152, n155, n158, n161, n164, n167, n170, n173, n176,
         n179, n182, n185, n188, n191, n194, n197, n200, n203, n206, n209,
         n212, n215, n218, n221, n224, n227, n230, n233, n236, n239, n242,
         n245, n248, n251, n254, n257, n260, n263, n266, n269, n272, n275,
         n278, n281, n285, n289, n291, n293, n295, n297, n299, n301, n303,
         n305, n307, n309, n311, n313, n315, n317, n319, n321, n323, n325,
         n327, n329, n331, n333, n335, n337, n339, n341, n343, n345, n347,
         n349, n351, n353, n355, n357, n359, n361, n363, n366, n369, n372,
         n375, n378, n381, n384, n387, n390, n393, n396, n399, n402, n405,
         n408, n411, n414, n417, n420, n423, n426, n429, n432, n435, n438,
         n441, n444, n447, n450, n453, n456, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n515, n517, n519, n521, n523, n525, n527, n529, n531, n533,
         n535, n537, n539, n541, n543, n545, n547, n549, n552, n555, n558,
         n561, n564, n567, n570, n573, n575, n578, n581, n584, n587, n590,
         n593, n596, n598, n600, n602, n605, n608, n611, n614, n617, n620,
         n622, n624, n626, n628, n630, n632, n634, n636, n638, n640, n642,
         n644, n646, n648, n650, n652, n654, n656, n658, n660, n662, n664,
         n666, n668, n670, n672, n674, n676, n678, n680, n682, n684, n686,
         n688, n690, n692, n694, n697, n700, n703, n706, n709, n712, n715,
         n718, n721, n724, n727, n730, n733, n736, n739, n742, n745, n748,
         n751, n754, n757, n760, n763, n766, n769, n772, n775, n778, n781,
         n784, n787, n790, n792, n794, n796, n798, n800, n802, n804, n806,
         n808, n810, n812, n814, n816, n818, n820, n822, n824, n826, n828,
         n830, n832, n834, n836, n838, n840, n842, n844, n846, n848, n850,
         n852, n854, n856, n858, n860, n862, n864, n866, n868, n870, n872,
         n874, n876, n878, n880, n883, n886, n889, n892, n895, n898, n901,
         n904, n906, n909, n912, n915, n918, n921, n924, n927, n929, n931,
         n935, n939, n941, n944, n947, n950, n953, n956, n959, n961, n963,
         n965, n967, n969, n971, n973, n975, n977, n979, n981, n983, n985,
         n987, n989, n991, n993, n995, n997, n999, n1001, n1003, n1005, n1007,
         n1009, n1011, n1013, n1015, n1017, n1019, n1021, n1023, n1025, n1027,
         n1029, n1031, n1033, n1036, n1039, n1042, n1045, n1048, n1051, n1054,
         n1057, n1060, n1063, n1066, n1069, n1072, n1075, n1078, n1081, n1084,
         n1087, n1090, n1093, n1096, n1099, n1102, n1105, n1108, n1111, n1114,
         n1117, n1120, n1123, n1126, n1129, n1131, n1133, n1135, n1137, n1139,
         n1141, n1143, n1145, n1147, n1149, n1151, n1153, n1155, n1157, n1159,
         n1161, n1163, n1165, n1167, n1169, n1171, n1173, n1175, n1177, n1179,
         n1181, n1183, n1185, n1187, n1189, n1191, n1193, n1195, n1197, n1199,
         n1201, n1203, n1205, n1207, n1209, n1211, n1213, n1215, n1217, n1219,
         n1222, n1225, n1228, n1231, n1234, n1237, n1240, n1243, n1245, n1248,
         n1251, n1254, n1257, n1260, n1263, n1266, n1268, n1270, n1274, n1278,
         n1280, n1283, n1286, n1289, n1292, n1295, n1298, n1300, n1302, n1304,
         n1306, n1308, n1310, n1312, n1314, n1316, n1318, n1320, n1322, n1324,
         n1326, n1328, n1330, n1332, n1334, n1336, n1338, n1340, n1342, n1344,
         n1346, n1348, n1350, n1352, n1354, n1356, n1358, n1360, n1362, n1364,
         n1366, n1368, n1370, n1372, n1374, n1376, n1378, n1380, n1382, n1384,
         n1386, n1388, n1390, n1392, n1394, n1396, n1398, n1400, n1402, n1404,
         n1406, n1408, n1410, n1412, n1414, n1416, n1418, n1420, n1422, n1424,
         n1426, n1428, n1430, n1432, n1434, n1436, n1438, n1440, n1442, n1444,
         n1446, n1448, n1450, n1452, n1454, n1456, n1458, n1460, n1462, n1464,
         n1466, n1468, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483;
  assign issueqPacket0_o_138 = renamedPacket0_i[138];
  assign issueqPacket0_o_131 = renamedPacket0_i[131];
  assign issueqPacket0_o_130 = renamedPacket0_i[130];
  assign issueqPacket0_o_122 = renamedPacket0_i[122];
  assign issueqPacket0_o_36 = renamedPacket0_i[36];
  assign issueqPacket0_o_35 = renamedPacket0_i[35];
  assign issueqPacket0_o_34 = renamedPacket0_i[34];
  assign issueqPacket0_o_33 = renamedPacket0_i[33];
  assign issueqPacket0_o_32 = renamedPacket0_i[32];
  assign issueqPacket0_o_31 = renamedPacket0_i[31];
  assign issueqPacket0_o_30 = renamedPacket0_i[30];
  assign issueqPacket0_o_29 = renamedPacket0_i[29];
  assign issueqPacket0_o_28 = renamedPacket0_i[28];
  assign issueqPacket0_o_27 = renamedPacket0_i[27];
  assign issueqPacket0_o_26 = renamedPacket0_i[26];
  assign issueqPacket0_o_25 = renamedPacket0_i[25];
  assign issueqPacket0_o_24 = renamedPacket0_i[24];
  assign issueqPacket0_o_23 = renamedPacket0_i[23];
  assign issueqPacket0_o_22 = renamedPacket0_i[22];
  assign issueqPacket0_o_21 = renamedPacket0_i[21];
  assign issueqPacket0_o_20 = renamedPacket0_i[20];
  assign issueqPacket0_o_19 = renamedPacket0_i[19];
  assign issueqPacket0_o_18 = renamedPacket0_i[18];
  assign issueqPacket0_o_17 = renamedPacket0_i[17];
  assign issueqPacket0_o_16 = renamedPacket0_i[16];
  assign issueqPacket0_o_15 = renamedPacket0_i[15];
  assign issueqPacket0_o_14 = renamedPacket0_i[14];
  assign issueqPacket0_o_13 = renamedPacket0_i[13];
  assign issueqPacket0_o_12 = renamedPacket0_i[12];
  assign issueqPacket0_o_11 = renamedPacket0_i[11];
  assign issueqPacket0_o_10 = renamedPacket0_i[10];
  assign issueqPacket0_o_9 = renamedPacket0_i[9];
  assign issueqPacket0_o_8 = renamedPacket0_i[8];
  assign issueqPacket0_o_7 = renamedPacket0_i[7];
  assign issueqPacket0_o_6 = renamedPacket0_i[6];
  assign issueqPacket0_o_5 = renamedPacket0_i[5];
  assign issueqPacket0_o_4 = renamedPacket0_i[4];
  assign issueqPacket0_o_3 = renamedPacket0_i[3];
  assign issueqPacket0_o_2 = renamedPacket0_i[2];
  assign issueqPacket0_o_1 = renamedPacket0_i[1];
  assign issueqPacket0_o_0 = renamedPacket0_i[0];
  assign issueqPacket1_o_144 = renamedPacket1_i[144];
  assign issueqPacket1_o_143 = renamedPacket1_i[143];
  assign issueqPacket1_o_142 = renamedPacket1_i[142];
  assign issueqPacket1_o_141 = renamedPacket1_i[141];
  assign issueqPacket1_o_140 = renamedPacket1_i[140];
  assign issueqPacket1_o_139 = renamedPacket1_i[139];
  assign issueqPacket1_o_138 = renamedPacket1_i[138];
  assign issueqPacket1_o_137 = renamedPacket1_i[137];
  assign issueqPacket1_o_136 = renamedPacket1_i[136];
  assign issueqPacket2_o_144 = renamedPacket2_i[144];
  assign issueqPacket2_o_143 = renamedPacket2_i[143];
  assign issueqPacket2_o_142 = renamedPacket2_i[142];
  assign issueqPacket2_o_141 = renamedPacket2_i[141];
  assign issueqPacket2_o_140 = renamedPacket2_i[140];
  assign issueqPacket2_o_139 = renamedPacket2_i[139];
  assign issueqPacket2_o_138 = renamedPacket2_i[138];
  assign issueqPacket2_o_137 = renamedPacket2_i[137];
  assign issueqPacket2_o_136 = renamedPacket2_i[136];
  assign issueqPacket3_o_144 = renamedPacket3_i[144];
  assign issueqPacket3_o_143 = renamedPacket3_i[143];
  assign issueqPacket3_o_142 = renamedPacket3_i[142];
  assign issueqPacket3_o_141 = renamedPacket3_i[141];
  assign issueqPacket3_o_140 = renamedPacket3_i[140];
  assign issueqPacket3_o_139 = renamedPacket3_i[139];
  assign issueqPacket3_o_138 = renamedPacket3_i[138];
  assign N44 = activeListCnt_i[1];
  assign N43 = activeListCnt_i[0];
  assign N37 = issueQueueCnt_i[1];
  assign N36 = issueQueueCnt_i[0];

  AND2X1 U28 ( .IN1(renamedPacket3_i[135]), .IN2(n61), .Q(lsqPacket3_o[5]) );
  AND2X1 U29 ( .IN1(renamedPacket3_i[134]), .IN2(n62), .Q(lsqPacket3_o[4]) );
  AND2X1 U30 ( .IN1(renamedPacket3_i[133]), .IN2(n63), .Q(lsqPacket3_o[3]) );
  AND2X1 U31 ( .IN1(renamedPacket3_i[132]), .IN2(n64), .Q(lsqPacket3_o[2]) );
  AND2X1 U32 ( .IN1(renamedPacket2_i[135]), .IN2(n61), .Q(lsqPacket2_o[5]) );
  AND2X1 U33 ( .IN1(renamedPacket2_i[134]), .IN2(n62), .Q(lsqPacket2_o[4]) );
  AND2X1 U34 ( .IN1(renamedPacket2_i[133]), .IN2(n63), .Q(lsqPacket2_o[3]) );
  AND2X1 U35 ( .IN1(renamedPacket2_i[132]), .IN2(n64), .Q(lsqPacket2_o[2]) );
  AND2X1 U36 ( .IN1(renamedPacket1_i[135]), .IN2(n61), .Q(lsqPacket1_o[5]) );
  AND2X1 U37 ( .IN1(renamedPacket1_i[134]), .IN2(n62), .Q(lsqPacket1_o[4]) );
  AND2X1 U38 ( .IN1(renamedPacket1_i[133]), .IN2(n63), .Q(lsqPacket1_o[3]) );
  AND2X1 U39 ( .IN1(renamedPacket1_i[132]), .IN2(n64), .Q(lsqPacket1_o[2]) );
  AND2X1 U40 ( .IN1(renamedPacket0_i[135]), .IN2(n61), .Q(lsqPacket0_o[5]) );
  NAND3X0 U41 ( .IN1(ctrlVerifiedSMTid_i[1]), .IN2(ctrlVerifiedSMTid_i[0]), 
        .IN3(ctrlVerified_i), .QN(n61) );
  AND2X1 U42 ( .IN1(renamedPacket0_i[134]), .IN2(n62), .Q(lsqPacket0_o[4]) );
  NAND3X0 U43 ( .IN1(ctrlVerifiedSMTid_i[1]), .IN2(n1479), .IN3(ctrlVerified_i), .QN(n62) );
  AND2X1 U44 ( .IN1(renamedPacket0_i[133]), .IN2(n63), .Q(lsqPacket0_o[3]) );
  NAND3X0 U45 ( .IN1(ctrlVerifiedSMTid_i[0]), .IN2(n1478), .IN3(ctrlVerified_i), .QN(n63) );
  AND2X1 U46 ( .IN1(renamedPacket0_i[132]), .IN2(n64), .Q(lsqPacket0_o[2]) );
  NAND3X0 U47 ( .IN1(n1479), .IN2(n1478), .IN3(ctrlVerified_i), .QN(n64) );
  AND2X1 U48 ( .IN1(n65), .IN2(renameReady_i), .Q(backEndReady_o) );
  OR4X1 U49 ( .IN1(stall1), .IN2(stall0), .IN3(stall3), .IN4(stall2), .Q(
        stallfrontEnd_o) );
  FADDX1 \add_288/U1_1  ( .A(loadQueueCnt_i[1]), .B(\loadCnt[1] ), .CI(
        \add_288/carry[1] ), .CO(\add_288/carry[2] ), .S(N23) );
  FADDX1 \add_288/U1_2  ( .A(loadQueueCnt_i[2]), .B(\loadCnt[2] ), .CI(
        \add_288/carry[2] ), .CO(\add_288/carry[3] ), .S(N24) );
  FADDX1 \add_289/U1_1  ( .A(storeQueueCnt_i[1]), .B(\storeCnt[1] ), .CI(
        \add_289/carry[1] ), .CO(\add_289/carry[2] ), .S(N30) );
  FADDX1 \add_289/U1_2  ( .A(storeQueueCnt_i[2]), .B(\storeCnt[2] ), .CI(
        \add_289/carry[2] ), .CO(\add_289/carry[3] ), .S(N31) );
  INVX0 U50 ( .INP(lsqPacket3_o[2]), .ZN(n66) );
  INVX0 U51 ( .INP(lsqPacket2_o[2]), .ZN(n78) );
  INVX0 U52 ( .INP(lsqPacket1_o[2]), .ZN(n90) );
  INVX0 U53 ( .INP(lsqPacket0_o[2]), .ZN(n102) );
  INVX0 U54 ( .INP(lsqPacket3_o[3]), .ZN(n69) );
  INVX0 U55 ( .INP(lsqPacket2_o[3]), .ZN(n81) );
  INVX0 U56 ( .INP(lsqPacket1_o[3]), .ZN(n93) );
  INVX0 U57 ( .INP(lsqPacket0_o[3]), .ZN(n105) );
  INVX0 U58 ( .INP(lsqPacket3_o[4]), .ZN(n72) );
  INVX0 U59 ( .INP(lsqPacket2_o[4]), .ZN(n84) );
  INVX0 U60 ( .INP(lsqPacket1_o[4]), .ZN(n96) );
  INVX0 U61 ( .INP(lsqPacket0_o[4]), .ZN(n108) );
  INVX0 U62 ( .INP(lsqPacket3_o[5]), .ZN(n75) );
  INVX0 U63 ( .INP(lsqPacket2_o[5]), .ZN(n87) );
  INVX0 U64 ( .INP(lsqPacket1_o[5]), .ZN(n99) );
  INVX0 U65 ( .INP(lsqPacket0_o[5]), .ZN(n111) );
  INVX0 U66 ( .INP(renamedPacket3_i[37]), .ZN(n363) );
  INVX0 U67 ( .INP(renamedPacket3_i[38]), .ZN(n366) );
  INVX0 U68 ( .INP(renamedPacket3_i[39]), .ZN(n369) );
  INVX0 U69 ( .INP(renamedPacket3_i[40]), .ZN(n372) );
  INVX0 U70 ( .INP(renamedPacket3_i[41]), .ZN(n375) );
  INVX0 U71 ( .INP(renamedPacket3_i[42]), .ZN(n378) );
  INVX0 U72 ( .INP(renamedPacket3_i[43]), .ZN(n381) );
  INVX0 U73 ( .INP(renamedPacket3_i[44]), .ZN(n384) );
  INVX0 U74 ( .INP(renamedPacket3_i[45]), .ZN(n387) );
  INVX0 U75 ( .INP(renamedPacket3_i[46]), .ZN(n390) );
  INVX0 U76 ( .INP(renamedPacket3_i[47]), .ZN(n393) );
  INVX0 U77 ( .INP(renamedPacket3_i[48]), .ZN(n396) );
  INVX0 U78 ( .INP(renamedPacket3_i[49]), .ZN(n399) );
  INVX0 U79 ( .INP(renamedPacket3_i[50]), .ZN(n402) );
  INVX0 U80 ( .INP(renamedPacket3_i[51]), .ZN(n405) );
  INVX0 U81 ( .INP(renamedPacket3_i[52]), .ZN(n408) );
  INVX0 U82 ( .INP(renamedPacket3_i[53]), .ZN(n411) );
  INVX0 U83 ( .INP(renamedPacket3_i[114]), .ZN(n549) );
  INVX0 U84 ( .INP(renamedPacket3_i[115]), .ZN(n552) );
  INVX0 U85 ( .INP(renamedPacket3_i[116]), .ZN(n555) );
  INVX0 U86 ( .INP(renamedPacket3_i[117]), .ZN(n558) );
  INVX0 U87 ( .INP(renamedPacket3_i[118]), .ZN(n561) );
  INVX0 U88 ( .INP(renamedPacket3_i[119]), .ZN(n564) );
  INVX0 U89 ( .INP(renamedPacket3_i[120]), .ZN(n567) );
  INVX0 U90 ( .INP(renamedPacket3_i[121]), .ZN(n570) );
  INVX0 U91 ( .INP(renamedPacket3_i[123]), .ZN(n575) );
  INVX0 U92 ( .INP(renamedPacket3_i[124]), .ZN(n578) );
  INVX0 U93 ( .INP(renamedPacket3_i[125]), .ZN(n581) );
  INVX0 U94 ( .INP(renamedPacket3_i[126]), .ZN(n584) );
  INVX0 U95 ( .INP(renamedPacket3_i[127]), .ZN(n587) );
  INVX0 U96 ( .INP(renamedPacket3_i[128]), .ZN(n590) );
  INVX0 U97 ( .INP(renamedPacket3_i[129]), .ZN(n593) );
  INVX0 U98 ( .INP(issueqPacket3_o_139), .ZN(n602) );
  INVX0 U99 ( .INP(issueqPacket3_o_140), .ZN(n605) );
  INVX0 U100 ( .INP(issueqPacket3_o_141), .ZN(n608) );
  INVX0 U101 ( .INP(issueqPacket3_o_142), .ZN(n611) );
  INVX0 U102 ( .INP(issueqPacket3_o_143), .ZN(n614) );
  INVX0 U103 ( .INP(issueqPacket3_o_144), .ZN(n617) );
  INVX0 U104 ( .INP(renamedPacket2_i[37]), .ZN(n694) );
  INVX0 U105 ( .INP(renamedPacket2_i[38]), .ZN(n697) );
  INVX0 U106 ( .INP(renamedPacket2_i[39]), .ZN(n700) );
  INVX0 U107 ( .INP(renamedPacket2_i[40]), .ZN(n703) );
  INVX0 U108 ( .INP(renamedPacket2_i[41]), .ZN(n706) );
  INVX0 U109 ( .INP(renamedPacket2_i[42]), .ZN(n709) );
  INVX0 U110 ( .INP(renamedPacket2_i[43]), .ZN(n712) );
  INVX0 U111 ( .INP(renamedPacket2_i[44]), .ZN(n715) );
  INVX0 U112 ( .INP(renamedPacket2_i[45]), .ZN(n718) );
  INVX0 U113 ( .INP(renamedPacket2_i[46]), .ZN(n721) );
  INVX0 U114 ( .INP(renamedPacket2_i[47]), .ZN(n724) );
  INVX0 U115 ( .INP(renamedPacket2_i[48]), .ZN(n727) );
  INVX0 U116 ( .INP(renamedPacket2_i[49]), .ZN(n730) );
  INVX0 U117 ( .INP(renamedPacket2_i[50]), .ZN(n733) );
  INVX0 U118 ( .INP(renamedPacket2_i[51]), .ZN(n736) );
  INVX0 U119 ( .INP(renamedPacket2_i[52]), .ZN(n739) );
  INVX0 U120 ( .INP(renamedPacket2_i[53]), .ZN(n742) );
  INVX0 U121 ( .INP(renamedPacket2_i[54]), .ZN(n745) );
  INVX0 U122 ( .INP(renamedPacket2_i[55]), .ZN(n748) );
  INVX0 U123 ( .INP(renamedPacket2_i[56]), .ZN(n751) );
  INVX0 U124 ( .INP(renamedPacket2_i[57]), .ZN(n754) );
  INVX0 U125 ( .INP(renamedPacket2_i[58]), .ZN(n757) );
  INVX0 U126 ( .INP(renamedPacket2_i[59]), .ZN(n760) );
  INVX0 U127 ( .INP(renamedPacket2_i[60]), .ZN(n763) );
  INVX0 U128 ( .INP(renamedPacket2_i[61]), .ZN(n766) );
  INVX0 U129 ( .INP(renamedPacket2_i[62]), .ZN(n769) );
  INVX0 U130 ( .INP(renamedPacket2_i[63]), .ZN(n772) );
  INVX0 U131 ( .INP(renamedPacket2_i[64]), .ZN(n775) );
  INVX0 U132 ( .INP(renamedPacket2_i[65]), .ZN(n778) );
  INVX0 U133 ( .INP(renamedPacket2_i[66]), .ZN(n781) );
  INVX0 U134 ( .INP(renamedPacket2_i[67]), .ZN(n784) );
  INVX0 U135 ( .INP(renamedPacket2_i[68]), .ZN(n787) );
  INVX0 U136 ( .INP(renamedPacket2_i[114]), .ZN(n880) );
  INVX0 U137 ( .INP(renamedPacket2_i[115]), .ZN(n883) );
  INVX0 U138 ( .INP(renamedPacket2_i[116]), .ZN(n886) );
  INVX0 U139 ( .INP(renamedPacket2_i[117]), .ZN(n889) );
  INVX0 U140 ( .INP(renamedPacket2_i[118]), .ZN(n892) );
  INVX0 U141 ( .INP(renamedPacket2_i[119]), .ZN(n895) );
  INVX0 U142 ( .INP(renamedPacket2_i[120]), .ZN(n898) );
  INVX0 U143 ( .INP(renamedPacket2_i[121]), .ZN(n901) );
  INVX0 U144 ( .INP(renamedPacket2_i[123]), .ZN(n906) );
  INVX0 U145 ( .INP(renamedPacket2_i[124]), .ZN(n909) );
  INVX0 U146 ( .INP(renamedPacket2_i[125]), .ZN(n912) );
  INVX0 U147 ( .INP(renamedPacket2_i[126]), .ZN(n915) );
  INVX0 U148 ( .INP(renamedPacket2_i[127]), .ZN(n918) );
  INVX0 U149 ( .INP(renamedPacket2_i[128]), .ZN(n921) );
  INVX0 U150 ( .INP(renamedPacket2_i[129]), .ZN(n924) );
  INVX0 U151 ( .INP(issueqPacket2_o_139), .ZN(n941) );
  INVX0 U152 ( .INP(issueqPacket2_o_140), .ZN(n944) );
  INVX0 U153 ( .INP(issueqPacket2_o_141), .ZN(n947) );
  INVX0 U154 ( .INP(issueqPacket2_o_142), .ZN(n950) );
  INVX0 U155 ( .INP(issueqPacket2_o_143), .ZN(n953) );
  INVX0 U156 ( .INP(issueqPacket2_o_144), .ZN(n956) );
  INVX0 U157 ( .INP(renamedPacket1_i[37]), .ZN(n1033) );
  INVX0 U158 ( .INP(renamedPacket1_i[38]), .ZN(n1036) );
  INVX0 U159 ( .INP(renamedPacket1_i[39]), .ZN(n1039) );
  INVX0 U160 ( .INP(renamedPacket1_i[40]), .ZN(n1042) );
  INVX0 U161 ( .INP(renamedPacket1_i[41]), .ZN(n1045) );
  INVX0 U162 ( .INP(renamedPacket1_i[42]), .ZN(n1048) );
  INVX0 U163 ( .INP(renamedPacket1_i[43]), .ZN(n1051) );
  INVX0 U164 ( .INP(renamedPacket1_i[44]), .ZN(n1054) );
  INVX0 U165 ( .INP(renamedPacket1_i[45]), .ZN(n1057) );
  INVX0 U166 ( .INP(renamedPacket1_i[46]), .ZN(n1060) );
  INVX0 U167 ( .INP(renamedPacket1_i[47]), .ZN(n1063) );
  INVX0 U168 ( .INP(renamedPacket1_i[48]), .ZN(n1066) );
  INVX0 U169 ( .INP(renamedPacket1_i[49]), .ZN(n1069) );
  INVX0 U170 ( .INP(renamedPacket1_i[50]), .ZN(n1072) );
  INVX0 U171 ( .INP(renamedPacket1_i[51]), .ZN(n1075) );
  INVX0 U172 ( .INP(renamedPacket1_i[52]), .ZN(n1078) );
  INVX0 U173 ( .INP(renamedPacket1_i[53]), .ZN(n1081) );
  INVX0 U174 ( .INP(renamedPacket1_i[54]), .ZN(n1084) );
  INVX0 U175 ( .INP(renamedPacket1_i[55]), .ZN(n1087) );
  INVX0 U176 ( .INP(renamedPacket1_i[56]), .ZN(n1090) );
  INVX0 U177 ( .INP(renamedPacket1_i[57]), .ZN(n1093) );
  INVX0 U178 ( .INP(renamedPacket1_i[58]), .ZN(n1096) );
  INVX0 U179 ( .INP(renamedPacket1_i[59]), .ZN(n1099) );
  INVX0 U180 ( .INP(renamedPacket1_i[60]), .ZN(n1102) );
  INVX0 U181 ( .INP(renamedPacket1_i[61]), .ZN(n1105) );
  INVX0 U182 ( .INP(renamedPacket1_i[62]), .ZN(n1108) );
  INVX0 U183 ( .INP(renamedPacket1_i[63]), .ZN(n1111) );
  INVX0 U184 ( .INP(renamedPacket1_i[64]), .ZN(n1114) );
  INVX0 U185 ( .INP(renamedPacket1_i[65]), .ZN(n1117) );
  INVX0 U186 ( .INP(renamedPacket1_i[66]), .ZN(n1120) );
  INVX0 U187 ( .INP(renamedPacket1_i[67]), .ZN(n1123) );
  INVX0 U188 ( .INP(renamedPacket1_i[68]), .ZN(n1126) );
  INVX0 U189 ( .INP(renamedPacket1_i[114]), .ZN(n1219) );
  INVX0 U190 ( .INP(renamedPacket1_i[115]), .ZN(n1222) );
  INVX0 U191 ( .INP(renamedPacket1_i[116]), .ZN(n1225) );
  INVX0 U192 ( .INP(renamedPacket1_i[117]), .ZN(n1228) );
  INVX0 U193 ( .INP(renamedPacket1_i[118]), .ZN(n1231) );
  INVX0 U194 ( .INP(renamedPacket1_i[119]), .ZN(n1234) );
  INVX0 U195 ( .INP(renamedPacket1_i[120]), .ZN(n1237) );
  INVX0 U196 ( .INP(renamedPacket1_i[121]), .ZN(n1240) );
  INVX0 U197 ( .INP(renamedPacket1_i[123]), .ZN(n1245) );
  INVX0 U198 ( .INP(renamedPacket1_i[124]), .ZN(n1248) );
  INVX0 U199 ( .INP(renamedPacket1_i[125]), .ZN(n1251) );
  INVX0 U200 ( .INP(renamedPacket1_i[126]), .ZN(n1254) );
  INVX0 U201 ( .INP(renamedPacket1_i[127]), .ZN(n1257) );
  INVX0 U202 ( .INP(renamedPacket1_i[128]), .ZN(n1260) );
  INVX0 U203 ( .INP(renamedPacket1_i[129]), .ZN(n1263) );
  INVX0 U204 ( .INP(issueqPacket1_o_139), .ZN(n1280) );
  INVX0 U205 ( .INP(issueqPacket1_o_140), .ZN(n1283) );
  INVX0 U206 ( .INP(issueqPacket1_o_141), .ZN(n1286) );
  INVX0 U207 ( .INP(issueqPacket1_o_142), .ZN(n1289) );
  INVX0 U208 ( .INP(issueqPacket1_o_143), .ZN(n1292) );
  INVX0 U209 ( .INP(issueqPacket1_o_144), .ZN(n1295) );
  INVX0 U210 ( .INP(renamedPacket0_i[37]), .ZN(n185) );
  INVX0 U211 ( .INP(renamedPacket0_i[38]), .ZN(n188) );
  INVX0 U212 ( .INP(renamedPacket0_i[39]), .ZN(n191) );
  INVX0 U213 ( .INP(renamedPacket0_i[40]), .ZN(n194) );
  INVX0 U214 ( .INP(renamedPacket0_i[41]), .ZN(n197) );
  INVX0 U215 ( .INP(renamedPacket0_i[42]), .ZN(n200) );
  INVX0 U216 ( .INP(renamedPacket0_i[43]), .ZN(n203) );
  INVX0 U217 ( .INP(renamedPacket0_i[44]), .ZN(n206) );
  INVX0 U218 ( .INP(renamedPacket0_i[45]), .ZN(n209) );
  INVX0 U219 ( .INP(renamedPacket0_i[46]), .ZN(n212) );
  INVX0 U220 ( .INP(renamedPacket0_i[47]), .ZN(n215) );
  INVX0 U221 ( .INP(renamedPacket0_i[48]), .ZN(n218) );
  INVX0 U222 ( .INP(renamedPacket0_i[49]), .ZN(n221) );
  INVX0 U223 ( .INP(renamedPacket0_i[50]), .ZN(n224) );
  INVX0 U224 ( .INP(renamedPacket0_i[51]), .ZN(n227) );
  INVX0 U225 ( .INP(renamedPacket0_i[52]), .ZN(n230) );
  INVX0 U226 ( .INP(renamedPacket0_i[53]), .ZN(n233) );
  INVX0 U227 ( .INP(renamedPacket0_i[54]), .ZN(n236) );
  INVX0 U228 ( .INP(renamedPacket0_i[55]), .ZN(n239) );
  INVX0 U229 ( .INP(renamedPacket0_i[56]), .ZN(n242) );
  INVX0 U230 ( .INP(renamedPacket0_i[57]), .ZN(n245) );
  INVX0 U231 ( .INP(renamedPacket0_i[58]), .ZN(n248) );
  INVX0 U232 ( .INP(renamedPacket0_i[59]), .ZN(n251) );
  INVX0 U233 ( .INP(renamedPacket0_i[60]), .ZN(n254) );
  INVX0 U234 ( .INP(renamedPacket0_i[61]), .ZN(n257) );
  INVX0 U235 ( .INP(renamedPacket0_i[62]), .ZN(n260) );
  INVX0 U236 ( .INP(renamedPacket0_i[63]), .ZN(n263) );
  INVX0 U237 ( .INP(renamedPacket0_i[64]), .ZN(n266) );
  INVX0 U238 ( .INP(renamedPacket0_i[65]), .ZN(n269) );
  INVX0 U239 ( .INP(renamedPacket0_i[66]), .ZN(n272) );
  INVX0 U240 ( .INP(renamedPacket0_i[67]), .ZN(n275) );
  INVX0 U241 ( .INP(renamedPacket0_i[68]), .ZN(n278) );
  INVX0 U242 ( .INP(renamedPacket0_i[114]), .ZN(n122) );
  INVX0 U243 ( .INP(renamedPacket0_i[115]), .ZN(n146) );
  INVX0 U244 ( .INP(renamedPacket0_i[116]), .ZN(n149) );
  INVX0 U245 ( .INP(renamedPacket0_i[117]), .ZN(n152) );
  INVX0 U246 ( .INP(renamedPacket0_i[118]), .ZN(n155) );
  INVX0 U247 ( .INP(renamedPacket0_i[119]), .ZN(n158) );
  INVX0 U248 ( .INP(renamedPacket0_i[120]), .ZN(n161) );
  INVX0 U249 ( .INP(renamedPacket0_i[121]), .ZN(n164) );
  INVX0 U250 ( .INP(renamedPacket0_i[123]), .ZN(n125) );
  INVX0 U251 ( .INP(renamedPacket0_i[124]), .ZN(n128) );
  INVX0 U252 ( .INP(renamedPacket0_i[125]), .ZN(n131) );
  INVX0 U253 ( .INP(renamedPacket0_i[126]), .ZN(n134) );
  INVX0 U254 ( .INP(renamedPacket0_i[127]), .ZN(n137) );
  INVX0 U255 ( .INP(renamedPacket0_i[128]), .ZN(n140) );
  INVX0 U256 ( .INP(renamedPacket0_i[129]), .ZN(n143) );
  INVX0 U257 ( .INP(renamedPacket0_i[139]), .ZN(n167) );
  INVX0 U258 ( .INP(renamedPacket0_i[140]), .ZN(n170) );
  INVX0 U259 ( .INP(renamedPacket0_i[141]), .ZN(n173) );
  INVX0 U260 ( .INP(renamedPacket0_i[142]), .ZN(n176) );
  INVX0 U261 ( .INP(renamedPacket0_i[143]), .ZN(n179) );
  INVX0 U262 ( .INP(renamedPacket0_i[144]), .ZN(n182) );
  INVX0 U263 ( .INP(renamedPacket3_i[136]), .ZN(n114) );
  INVX0 U264 ( .INP(renamedPacket3_i[137]), .ZN(n118) );
  INVX0 U265 ( .INP(issueqPacket2_o_136), .ZN(n931) );
  INVX0 U266 ( .INP(issueqPacket2_o_137), .ZN(n935) );
  INVX0 U267 ( .INP(issueqPacket1_o_136), .ZN(n1270) );
  INVX0 U268 ( .INP(issueqPacket1_o_137), .ZN(n1274) );
  INVX0 U269 ( .INP(renamedPacket0_i[136]), .ZN(n285) );
  INVX0 U270 ( .INP(renamedPacket0_i[137]), .ZN(n281) );
  INVX0 U271 ( .INP(n66), .ZN(updatedBranchMask3_o[0]) );
  INVX0 U272 ( .INP(n69), .ZN(updatedBranchMask3_o[1]) );
  INVX0 U273 ( .INP(n72), .ZN(updatedBranchMask3_o[2]) );
  INVX0 U274 ( .INP(n75), .ZN(updatedBranchMask3_o[3]) );
  INVX0 U275 ( .INP(n78), .ZN(updatedBranchMask2_o[0]) );
  INVX0 U276 ( .INP(n81), .ZN(updatedBranchMask2_o[1]) );
  INVX0 U277 ( .INP(n84), .ZN(updatedBranchMask2_o[2]) );
  INVX0 U278 ( .INP(n87), .ZN(updatedBranchMask2_o[3]) );
  INVX0 U279 ( .INP(n90), .ZN(updatedBranchMask1_o[0]) );
  INVX0 U280 ( .INP(n93), .ZN(updatedBranchMask1_o[1]) );
  INVX0 U281 ( .INP(n96), .ZN(updatedBranchMask1_o[2]) );
  INVX0 U282 ( .INP(n99), .ZN(updatedBranchMask1_o[3]) );
  INVX0 U283 ( .INP(n102), .ZN(updatedBranchMask0_o[0]) );
  INVX0 U284 ( .INP(n105), .ZN(updatedBranchMask0_o[1]) );
  INVX0 U285 ( .INP(n108), .ZN(updatedBranchMask0_o[2]) );
  INVX0 U286 ( .INP(n111), .ZN(updatedBranchMask0_o[3]) );
  INVX0 U287 ( .INP(n66), .ZN(issueqPacket3_o[132]) );
  INVX0 U288 ( .INP(n69), .ZN(issueqPacket3_o[133]) );
  INVX0 U289 ( .INP(n72), .ZN(issueqPacket3_o[134]) );
  INVX0 U290 ( .INP(n75), .ZN(issueqPacket3_o[135]) );
  INVX0 U291 ( .INP(n78), .ZN(issueqPacket2_o[132]) );
  INVX0 U292 ( .INP(n81), .ZN(issueqPacket2_o[133]) );
  INVX0 U293 ( .INP(n84), .ZN(issueqPacket2_o[134]) );
  INVX0 U294 ( .INP(n87), .ZN(issueqPacket2_o[135]) );
  INVX0 U295 ( .INP(n90), .ZN(issueqPacket1_o[132]) );
  INVX0 U296 ( .INP(n93), .ZN(issueqPacket1_o[133]) );
  INVX0 U297 ( .INP(n96), .ZN(issueqPacket1_o[134]) );
  INVX0 U298 ( .INP(n99), .ZN(issueqPacket1_o[135]) );
  INVX0 U299 ( .INP(n102), .ZN(issueqPacket0_o[132]) );
  INVX0 U300 ( .INP(n105), .ZN(issueqPacket0_o[133]) );
  INVX0 U301 ( .INP(n108), .ZN(issueqPacket0_o[134]) );
  INVX0 U302 ( .INP(n111), .ZN(issueqPacket0_o[135]) );
  INVX0 U303 ( .INP(n285), .ZN(lsqPacket0_o[0]) );
  INVX0 U304 ( .INP(n281), .ZN(lsqPacket0_o[1]) );
  INVX0 U305 ( .INP(n281), .ZN(alPacket0_o[53]) );
  INVX0 U306 ( .INP(n285), .ZN(alPacket0_o[54]) );
  INVX0 U307 ( .INP(n285), .ZN(issueqPacket0_o[136]) );
  INVX0 U308 ( .INP(n281), .ZN(issueqPacket0_o[137]) );
  INVX0 U309 ( .INP(n114), .ZN(lsqPacket3_o[0]) );
  INVX0 U310 ( .INP(n118), .ZN(lsqPacket3_o[1]) );
  INVX0 U311 ( .INP(n931), .ZN(lsqPacket2_o[0]) );
  INVX0 U312 ( .INP(n935), .ZN(lsqPacket2_o[1]) );
  INVX0 U313 ( .INP(n1270), .ZN(lsqPacket1_o[0]) );
  INVX0 U314 ( .INP(n1274), .ZN(lsqPacket1_o[1]) );
  INVX0 U315 ( .INP(n118), .ZN(alPacket3_o[53]) );
  INVX0 U316 ( .INP(n114), .ZN(alPacket3_o[54]) );
  INVX0 U317 ( .INP(n935), .ZN(alPacket2_o[53]) );
  INVX0 U318 ( .INP(n931), .ZN(alPacket2_o[54]) );
  INVX0 U319 ( .INP(n1274), .ZN(alPacket1_o[53]) );
  INVX0 U320 ( .INP(n1270), .ZN(alPacket1_o[54]) );
  INVX0 U321 ( .INP(n114), .ZN(issueqPacket3_o[136]) );
  INVX0 U322 ( .INP(n118), .ZN(issueqPacket3_o[137]) );
  INVX0 U323 ( .INP(n931), .ZN(issueqPacket2_o[136]) );
  INVX0 U324 ( .INP(n935), .ZN(issueqPacket2_o[137]) );
  INVX0 U325 ( .INP(n1270), .ZN(issueqPacket1_o[136]) );
  INVX0 U326 ( .INP(n1274), .ZN(issueqPacket1_o[137]) );
  INVX0 U327 ( .INP(n549), .ZN(alPacket3_o[0]) );
  INVX0 U328 ( .INP(n575), .ZN(alPacket3_o[1]) );
  INVX0 U329 ( .INP(n578), .ZN(alPacket3_o[2]) );
  INVX0 U330 ( .INP(n581), .ZN(alPacket3_o[3]) );
  INVX0 U331 ( .INP(n584), .ZN(alPacket3_o[4]) );
  INVX0 U332 ( .INP(n587), .ZN(alPacket3_o[5]) );
  INVX0 U333 ( .INP(n590), .ZN(alPacket3_o[6]) );
  INVX0 U334 ( .INP(n593), .ZN(alPacket3_o[7]) );
  INVX0 U335 ( .INP(n552), .ZN(alPacket3_o[8]) );
  INVX0 U336 ( .INP(n555), .ZN(alPacket3_o[9]) );
  INVX0 U337 ( .INP(n558), .ZN(alPacket3_o[10]) );
  INVX0 U338 ( .INP(n561), .ZN(alPacket3_o[11]) );
  INVX0 U339 ( .INP(n564), .ZN(alPacket3_o[12]) );
  INVX0 U340 ( .INP(n567), .ZN(alPacket3_o[13]) );
  INVX0 U341 ( .INP(n570), .ZN(alPacket3_o[14]) );
  INVX0 U342 ( .INP(n602), .ZN(alPacket3_o[15]) );
  INVX0 U343 ( .INP(n605), .ZN(alPacket3_o[16]) );
  INVX0 U344 ( .INP(n608), .ZN(alPacket3_o[17]) );
  INVX0 U345 ( .INP(n611), .ZN(alPacket3_o[18]) );
  INVX0 U346 ( .INP(n614), .ZN(alPacket3_o[19]) );
  INVX0 U347 ( .INP(n617), .ZN(alPacket3_o[20]) );
  INVX0 U348 ( .INP(n363), .ZN(alPacket3_o[21]) );
  INVX0 U349 ( .INP(n366), .ZN(alPacket3_o[22]) );
  INVX0 U350 ( .INP(n369), .ZN(alPacket3_o[23]) );
  INVX0 U351 ( .INP(n372), .ZN(alPacket3_o[24]) );
  INVX0 U352 ( .INP(n375), .ZN(alPacket3_o[25]) );
  INVX0 U353 ( .INP(n378), .ZN(alPacket3_o[26]) );
  INVX0 U354 ( .INP(n381), .ZN(alPacket3_o[27]) );
  INVX0 U355 ( .INP(n384), .ZN(alPacket3_o[28]) );
  INVX0 U356 ( .INP(n387), .ZN(alPacket3_o[29]) );
  INVX0 U357 ( .INP(n390), .ZN(alPacket3_o[30]) );
  INVX0 U358 ( .INP(n393), .ZN(alPacket3_o[31]) );
  INVX0 U359 ( .INP(n396), .ZN(alPacket3_o[32]) );
  INVX0 U360 ( .INP(n399), .ZN(alPacket3_o[33]) );
  INVX0 U361 ( .INP(n402), .ZN(alPacket3_o[34]) );
  INVX0 U362 ( .INP(n405), .ZN(alPacket3_o[35]) );
  INVX0 U363 ( .INP(n408), .ZN(alPacket3_o[36]) );
  INVX0 U364 ( .INP(n411), .ZN(alPacket3_o[37]) );
  INVX0 U365 ( .INP(n880), .ZN(alPacket2_o[0]) );
  INVX0 U366 ( .INP(n906), .ZN(alPacket2_o[1]) );
  INVX0 U367 ( .INP(n909), .ZN(alPacket2_o[2]) );
  INVX0 U368 ( .INP(n912), .ZN(alPacket2_o[3]) );
  INVX0 U369 ( .INP(n915), .ZN(alPacket2_o[4]) );
  INVX0 U370 ( .INP(n918), .ZN(alPacket2_o[5]) );
  INVX0 U371 ( .INP(n921), .ZN(alPacket2_o[6]) );
  INVX0 U372 ( .INP(n924), .ZN(alPacket2_o[7]) );
  INVX0 U373 ( .INP(n883), .ZN(alPacket2_o[8]) );
  INVX0 U374 ( .INP(n886), .ZN(alPacket2_o[9]) );
  INVX0 U375 ( .INP(n889), .ZN(alPacket2_o[10]) );
  INVX0 U376 ( .INP(n892), .ZN(alPacket2_o[11]) );
  INVX0 U377 ( .INP(n895), .ZN(alPacket2_o[12]) );
  INVX0 U378 ( .INP(n898), .ZN(alPacket2_o[13]) );
  INVX0 U379 ( .INP(n901), .ZN(alPacket2_o[14]) );
  INVX0 U380 ( .INP(n941), .ZN(alPacket2_o[15]) );
  INVX0 U381 ( .INP(n944), .ZN(alPacket2_o[16]) );
  INVX0 U382 ( .INP(n947), .ZN(alPacket2_o[17]) );
  INVX0 U383 ( .INP(n950), .ZN(alPacket2_o[18]) );
  INVX0 U384 ( .INP(n953), .ZN(alPacket2_o[19]) );
  INVX0 U385 ( .INP(n956), .ZN(alPacket2_o[20]) );
  INVX0 U386 ( .INP(n694), .ZN(alPacket2_o[21]) );
  INVX0 U387 ( .INP(n697), .ZN(alPacket2_o[22]) );
  INVX0 U388 ( .INP(n700), .ZN(alPacket2_o[23]) );
  INVX0 U389 ( .INP(n703), .ZN(alPacket2_o[24]) );
  INVX0 U390 ( .INP(n706), .ZN(alPacket2_o[25]) );
  INVX0 U391 ( .INP(n709), .ZN(alPacket2_o[26]) );
  INVX0 U392 ( .INP(n712), .ZN(alPacket2_o[27]) );
  INVX0 U393 ( .INP(n715), .ZN(alPacket2_o[28]) );
  INVX0 U394 ( .INP(n718), .ZN(alPacket2_o[29]) );
  INVX0 U395 ( .INP(n721), .ZN(alPacket2_o[30]) );
  INVX0 U396 ( .INP(n724), .ZN(alPacket2_o[31]) );
  INVX0 U397 ( .INP(n727), .ZN(alPacket2_o[32]) );
  INVX0 U398 ( .INP(n730), .ZN(alPacket2_o[33]) );
  INVX0 U399 ( .INP(n733), .ZN(alPacket2_o[34]) );
  INVX0 U400 ( .INP(n736), .ZN(alPacket2_o[35]) );
  INVX0 U401 ( .INP(n739), .ZN(alPacket2_o[36]) );
  INVX0 U402 ( .INP(n742), .ZN(alPacket2_o[37]) );
  INVX0 U403 ( .INP(n745), .ZN(alPacket2_o[38]) );
  INVX0 U404 ( .INP(n748), .ZN(alPacket2_o[39]) );
  INVX0 U405 ( .INP(n751), .ZN(alPacket2_o[40]) );
  INVX0 U406 ( .INP(n754), .ZN(alPacket2_o[41]) );
  INVX0 U407 ( .INP(n757), .ZN(alPacket2_o[42]) );
  INVX0 U408 ( .INP(n760), .ZN(alPacket2_o[43]) );
  INVX0 U409 ( .INP(n763), .ZN(alPacket2_o[44]) );
  INVX0 U410 ( .INP(n766), .ZN(alPacket2_o[45]) );
  INVX0 U411 ( .INP(n769), .ZN(alPacket2_o[46]) );
  INVX0 U412 ( .INP(n772), .ZN(alPacket2_o[47]) );
  INVX0 U413 ( .INP(n775), .ZN(alPacket2_o[48]) );
  INVX0 U414 ( .INP(n778), .ZN(alPacket2_o[49]) );
  INVX0 U415 ( .INP(n781), .ZN(alPacket2_o[50]) );
  INVX0 U416 ( .INP(n784), .ZN(alPacket2_o[51]) );
  INVX0 U417 ( .INP(n787), .ZN(alPacket2_o[52]) );
  INVX0 U418 ( .INP(n1219), .ZN(alPacket1_o[0]) );
  INVX0 U419 ( .INP(n1245), .ZN(alPacket1_o[1]) );
  INVX0 U420 ( .INP(n1248), .ZN(alPacket1_o[2]) );
  INVX0 U421 ( .INP(n1251), .ZN(alPacket1_o[3]) );
  INVX0 U422 ( .INP(n1254), .ZN(alPacket1_o[4]) );
  INVX0 U423 ( .INP(n1257), .ZN(alPacket1_o[5]) );
  INVX0 U424 ( .INP(n1260), .ZN(alPacket1_o[6]) );
  INVX0 U425 ( .INP(n1263), .ZN(alPacket1_o[7]) );
  INVX0 U426 ( .INP(n1222), .ZN(alPacket1_o[8]) );
  INVX0 U427 ( .INP(n1225), .ZN(alPacket1_o[9]) );
  INVX0 U428 ( .INP(n1228), .ZN(alPacket1_o[10]) );
  INVX0 U429 ( .INP(n1231), .ZN(alPacket1_o[11]) );
  INVX0 U430 ( .INP(n1234), .ZN(alPacket1_o[12]) );
  INVX0 U431 ( .INP(n1237), .ZN(alPacket1_o[13]) );
  INVX0 U432 ( .INP(n1240), .ZN(alPacket1_o[14]) );
  INVX0 U433 ( .INP(n1280), .ZN(alPacket1_o[15]) );
  INVX0 U434 ( .INP(n1283), .ZN(alPacket1_o[16]) );
  INVX0 U435 ( .INP(n1286), .ZN(alPacket1_o[17]) );
  INVX0 U436 ( .INP(n1289), .ZN(alPacket1_o[18]) );
  INVX0 U437 ( .INP(n1292), .ZN(alPacket1_o[19]) );
  INVX0 U438 ( .INP(n1295), .ZN(alPacket1_o[20]) );
  INVX0 U439 ( .INP(n1033), .ZN(alPacket1_o[21]) );
  INVX0 U440 ( .INP(n1036), .ZN(alPacket1_o[22]) );
  INVX0 U441 ( .INP(n1039), .ZN(alPacket1_o[23]) );
  INVX0 U442 ( .INP(n1042), .ZN(alPacket1_o[24]) );
  INVX0 U443 ( .INP(n1045), .ZN(alPacket1_o[25]) );
  INVX0 U444 ( .INP(n1048), .ZN(alPacket1_o[26]) );
  INVX0 U445 ( .INP(n1051), .ZN(alPacket1_o[27]) );
  INVX0 U446 ( .INP(n1054), .ZN(alPacket1_o[28]) );
  INVX0 U447 ( .INP(n1057), .ZN(alPacket1_o[29]) );
  INVX0 U448 ( .INP(n1060), .ZN(alPacket1_o[30]) );
  INVX0 U449 ( .INP(n1063), .ZN(alPacket1_o[31]) );
  INVX0 U450 ( .INP(n1066), .ZN(alPacket1_o[32]) );
  INVX0 U451 ( .INP(n1069), .ZN(alPacket1_o[33]) );
  INVX0 U452 ( .INP(n1072), .ZN(alPacket1_o[34]) );
  INVX0 U453 ( .INP(n1075), .ZN(alPacket1_o[35]) );
  INVX0 U454 ( .INP(n1078), .ZN(alPacket1_o[36]) );
  INVX0 U455 ( .INP(n1081), .ZN(alPacket1_o[37]) );
  INVX0 U456 ( .INP(n1084), .ZN(alPacket1_o[38]) );
  INVX0 U457 ( .INP(n1087), .ZN(alPacket1_o[39]) );
  INVX0 U458 ( .INP(n1090), .ZN(alPacket1_o[40]) );
  INVX0 U459 ( .INP(n1093), .ZN(alPacket1_o[41]) );
  INVX0 U460 ( .INP(n1096), .ZN(alPacket1_o[42]) );
  INVX0 U461 ( .INP(n1099), .ZN(alPacket1_o[43]) );
  INVX0 U462 ( .INP(n1102), .ZN(alPacket1_o[44]) );
  INVX0 U463 ( .INP(n1105), .ZN(alPacket1_o[45]) );
  INVX0 U464 ( .INP(n1108), .ZN(alPacket1_o[46]) );
  INVX0 U465 ( .INP(n1111), .ZN(alPacket1_o[47]) );
  INVX0 U466 ( .INP(n1114), .ZN(alPacket1_o[48]) );
  INVX0 U467 ( .INP(n1117), .ZN(alPacket1_o[49]) );
  INVX0 U468 ( .INP(n1120), .ZN(alPacket1_o[50]) );
  INVX0 U469 ( .INP(n1123), .ZN(alPacket1_o[51]) );
  INVX0 U470 ( .INP(n1126), .ZN(alPacket1_o[52]) );
  INVX0 U471 ( .INP(n122), .ZN(alPacket0_o[0]) );
  INVX0 U472 ( .INP(n125), .ZN(alPacket0_o[1]) );
  INVX0 U473 ( .INP(n128), .ZN(alPacket0_o[2]) );
  INVX0 U474 ( .INP(n131), .ZN(alPacket0_o[3]) );
  INVX0 U475 ( .INP(n134), .ZN(alPacket0_o[4]) );
  INVX0 U476 ( .INP(n137), .ZN(alPacket0_o[5]) );
  INVX0 U477 ( .INP(n140), .ZN(alPacket0_o[6]) );
  INVX0 U478 ( .INP(n143), .ZN(alPacket0_o[7]) );
  INVX0 U479 ( .INP(n146), .ZN(alPacket0_o[8]) );
  INVX0 U480 ( .INP(n149), .ZN(alPacket0_o[9]) );
  INVX0 U481 ( .INP(n152), .ZN(alPacket0_o[10]) );
  INVX0 U482 ( .INP(n155), .ZN(alPacket0_o[11]) );
  INVX0 U483 ( .INP(n158), .ZN(alPacket0_o[12]) );
  INVX0 U484 ( .INP(n161), .ZN(alPacket0_o[13]) );
  INVX0 U485 ( .INP(n164), .ZN(alPacket0_o[14]) );
  INVX0 U486 ( .INP(n167), .ZN(alPacket0_o[15]) );
  INVX0 U487 ( .INP(n170), .ZN(alPacket0_o[16]) );
  INVX0 U488 ( .INP(n173), .ZN(alPacket0_o[17]) );
  INVX0 U489 ( .INP(n176), .ZN(alPacket0_o[18]) );
  INVX0 U490 ( .INP(n179), .ZN(alPacket0_o[19]) );
  INVX0 U491 ( .INP(n182), .ZN(alPacket0_o[20]) );
  INVX0 U492 ( .INP(n185), .ZN(alPacket0_o[21]) );
  INVX0 U493 ( .INP(n188), .ZN(alPacket0_o[22]) );
  INVX0 U494 ( .INP(n191), .ZN(alPacket0_o[23]) );
  INVX0 U495 ( .INP(n194), .ZN(alPacket0_o[24]) );
  INVX0 U496 ( .INP(n197), .ZN(alPacket0_o[25]) );
  INVX0 U497 ( .INP(n200), .ZN(alPacket0_o[26]) );
  INVX0 U498 ( .INP(n203), .ZN(alPacket0_o[27]) );
  INVX0 U499 ( .INP(n206), .ZN(alPacket0_o[28]) );
  INVX0 U500 ( .INP(n209), .ZN(alPacket0_o[29]) );
  INVX0 U501 ( .INP(n212), .ZN(alPacket0_o[30]) );
  INVX0 U502 ( .INP(n215), .ZN(alPacket0_o[31]) );
  INVX0 U503 ( .INP(n218), .ZN(alPacket0_o[32]) );
  INVX0 U504 ( .INP(n221), .ZN(alPacket0_o[33]) );
  INVX0 U505 ( .INP(n224), .ZN(alPacket0_o[34]) );
  INVX0 U506 ( .INP(n227), .ZN(alPacket0_o[35]) );
  INVX0 U507 ( .INP(n230), .ZN(alPacket0_o[36]) );
  INVX0 U508 ( .INP(n233), .ZN(alPacket0_o[37]) );
  INVX0 U509 ( .INP(n236), .ZN(alPacket0_o[38]) );
  INVX0 U510 ( .INP(n239), .ZN(alPacket0_o[39]) );
  INVX0 U511 ( .INP(n242), .ZN(alPacket0_o[40]) );
  INVX0 U512 ( .INP(n245), .ZN(alPacket0_o[41]) );
  INVX0 U513 ( .INP(n248), .ZN(alPacket0_o[42]) );
  INVX0 U514 ( .INP(n251), .ZN(alPacket0_o[43]) );
  INVX0 U515 ( .INP(n254), .ZN(alPacket0_o[44]) );
  INVX0 U516 ( .INP(n257), .ZN(alPacket0_o[45]) );
  INVX0 U517 ( .INP(n260), .ZN(alPacket0_o[46]) );
  INVX0 U518 ( .INP(n263), .ZN(alPacket0_o[47]) );
  INVX0 U519 ( .INP(n266), .ZN(alPacket0_o[48]) );
  INVX0 U520 ( .INP(n269), .ZN(alPacket0_o[49]) );
  INVX0 U521 ( .INP(n272), .ZN(alPacket0_o[50]) );
  INVX0 U522 ( .INP(n275), .ZN(alPacket0_o[51]) );
  INVX0 U523 ( .INP(n278), .ZN(alPacket0_o[52]) );
  INVX0 U524 ( .INP(n363), .ZN(issueqPacket3_o[37]) );
  INVX0 U525 ( .INP(n366), .ZN(issueqPacket3_o[38]) );
  INVX0 U526 ( .INP(n369), .ZN(issueqPacket3_o[39]) );
  INVX0 U527 ( .INP(n372), .ZN(issueqPacket3_o[40]) );
  INVX0 U528 ( .INP(n375), .ZN(issueqPacket3_o[41]) );
  INVX0 U529 ( .INP(n378), .ZN(issueqPacket3_o[42]) );
  INVX0 U530 ( .INP(n381), .ZN(issueqPacket3_o[43]) );
  INVX0 U531 ( .INP(n384), .ZN(issueqPacket3_o[44]) );
  INVX0 U532 ( .INP(n387), .ZN(issueqPacket3_o[45]) );
  INVX0 U533 ( .INP(n390), .ZN(issueqPacket3_o[46]) );
  INVX0 U534 ( .INP(n393), .ZN(issueqPacket3_o[47]) );
  INVX0 U535 ( .INP(n396), .ZN(issueqPacket3_o[48]) );
  INVX0 U536 ( .INP(n399), .ZN(issueqPacket3_o[49]) );
  INVX0 U537 ( .INP(n402), .ZN(issueqPacket3_o[50]) );
  INVX0 U538 ( .INP(n405), .ZN(issueqPacket3_o[51]) );
  INVX0 U539 ( .INP(n408), .ZN(issueqPacket3_o[52]) );
  INVX0 U540 ( .INP(n411), .ZN(issueqPacket3_o[53]) );
  INVX0 U541 ( .INP(n549), .ZN(issueqPacket3_o[114]) );
  INVX0 U542 ( .INP(n552), .ZN(issueqPacket3_o[115]) );
  INVX0 U543 ( .INP(n555), .ZN(issueqPacket3_o[116]) );
  INVX0 U544 ( .INP(n558), .ZN(issueqPacket3_o[117]) );
  INVX0 U545 ( .INP(n561), .ZN(issueqPacket3_o[118]) );
  INVX0 U546 ( .INP(n564), .ZN(issueqPacket3_o[119]) );
  INVX0 U547 ( .INP(n567), .ZN(issueqPacket3_o[120]) );
  INVX0 U548 ( .INP(n570), .ZN(issueqPacket3_o[121]) );
  INVX0 U549 ( .INP(n575), .ZN(issueqPacket3_o[123]) );
  INVX0 U550 ( .INP(n578), .ZN(issueqPacket3_o[124]) );
  INVX0 U551 ( .INP(n581), .ZN(issueqPacket3_o[125]) );
  INVX0 U552 ( .INP(n584), .ZN(issueqPacket3_o[126]) );
  INVX0 U553 ( .INP(n587), .ZN(issueqPacket3_o[127]) );
  INVX0 U554 ( .INP(n590), .ZN(issueqPacket3_o[128]) );
  INVX0 U555 ( .INP(n593), .ZN(issueqPacket3_o[129]) );
  INVX0 U556 ( .INP(n602), .ZN(issueqPacket3_o[139]) );
  INVX0 U557 ( .INP(n605), .ZN(issueqPacket3_o[140]) );
  INVX0 U558 ( .INP(n608), .ZN(issueqPacket3_o[141]) );
  INVX0 U559 ( .INP(n611), .ZN(issueqPacket3_o[142]) );
  INVX0 U560 ( .INP(n614), .ZN(issueqPacket3_o[143]) );
  INVX0 U561 ( .INP(n617), .ZN(issueqPacket3_o[144]) );
  INVX0 U562 ( .INP(n694), .ZN(issueqPacket2_o[37]) );
  INVX0 U563 ( .INP(n697), .ZN(issueqPacket2_o[38]) );
  INVX0 U564 ( .INP(n700), .ZN(issueqPacket2_o[39]) );
  INVX0 U565 ( .INP(n703), .ZN(issueqPacket2_o[40]) );
  INVX0 U566 ( .INP(n706), .ZN(issueqPacket2_o[41]) );
  INVX0 U567 ( .INP(n709), .ZN(issueqPacket2_o[42]) );
  INVX0 U568 ( .INP(n712), .ZN(issueqPacket2_o[43]) );
  INVX0 U569 ( .INP(n715), .ZN(issueqPacket2_o[44]) );
  INVX0 U570 ( .INP(n718), .ZN(issueqPacket2_o[45]) );
  INVX0 U571 ( .INP(n721), .ZN(issueqPacket2_o[46]) );
  INVX0 U572 ( .INP(n724), .ZN(issueqPacket2_o[47]) );
  INVX0 U573 ( .INP(n727), .ZN(issueqPacket2_o[48]) );
  INVX0 U574 ( .INP(n730), .ZN(issueqPacket2_o[49]) );
  INVX0 U575 ( .INP(n733), .ZN(issueqPacket2_o[50]) );
  INVX0 U576 ( .INP(n736), .ZN(issueqPacket2_o[51]) );
  INVX0 U577 ( .INP(n739), .ZN(issueqPacket2_o[52]) );
  INVX0 U578 ( .INP(n742), .ZN(issueqPacket2_o[53]) );
  INVX0 U579 ( .INP(n745), .ZN(issueqPacket2_o[54]) );
  INVX0 U580 ( .INP(n748), .ZN(issueqPacket2_o[55]) );
  INVX0 U581 ( .INP(n751), .ZN(issueqPacket2_o[56]) );
  INVX0 U582 ( .INP(n754), .ZN(issueqPacket2_o[57]) );
  INVX0 U583 ( .INP(n757), .ZN(issueqPacket2_o[58]) );
  INVX0 U584 ( .INP(n760), .ZN(issueqPacket2_o[59]) );
  INVX0 U585 ( .INP(n763), .ZN(issueqPacket2_o[60]) );
  INVX0 U586 ( .INP(n766), .ZN(issueqPacket2_o[61]) );
  INVX0 U587 ( .INP(n769), .ZN(issueqPacket2_o[62]) );
  INVX0 U588 ( .INP(n772), .ZN(issueqPacket2_o[63]) );
  INVX0 U589 ( .INP(n775), .ZN(issueqPacket2_o[64]) );
  INVX0 U590 ( .INP(n778), .ZN(issueqPacket2_o[65]) );
  INVX0 U591 ( .INP(n781), .ZN(issueqPacket2_o[66]) );
  INVX0 U592 ( .INP(n784), .ZN(issueqPacket2_o[67]) );
  INVX0 U593 ( .INP(n787), .ZN(issueqPacket2_o[68]) );
  INVX0 U594 ( .INP(n880), .ZN(issueqPacket2_o[114]) );
  INVX0 U595 ( .INP(n883), .ZN(issueqPacket2_o[115]) );
  INVX0 U596 ( .INP(n886), .ZN(issueqPacket2_o[116]) );
  INVX0 U597 ( .INP(n889), .ZN(issueqPacket2_o[117]) );
  INVX0 U598 ( .INP(n892), .ZN(issueqPacket2_o[118]) );
  INVX0 U599 ( .INP(n895), .ZN(issueqPacket2_o[119]) );
  INVX0 U600 ( .INP(n898), .ZN(issueqPacket2_o[120]) );
  INVX0 U601 ( .INP(n901), .ZN(issueqPacket2_o[121]) );
  INVX0 U602 ( .INP(n906), .ZN(issueqPacket2_o[123]) );
  INVX0 U603 ( .INP(n909), .ZN(issueqPacket2_o[124]) );
  INVX0 U604 ( .INP(n912), .ZN(issueqPacket2_o[125]) );
  INVX0 U605 ( .INP(n915), .ZN(issueqPacket2_o[126]) );
  INVX0 U606 ( .INP(n918), .ZN(issueqPacket2_o[127]) );
  INVX0 U607 ( .INP(n921), .ZN(issueqPacket2_o[128]) );
  INVX0 U608 ( .INP(n924), .ZN(issueqPacket2_o[129]) );
  INVX0 U609 ( .INP(n941), .ZN(issueqPacket2_o[139]) );
  INVX0 U610 ( .INP(n944), .ZN(issueqPacket2_o[140]) );
  INVX0 U611 ( .INP(n947), .ZN(issueqPacket2_o[141]) );
  INVX0 U612 ( .INP(n950), .ZN(issueqPacket2_o[142]) );
  INVX0 U613 ( .INP(n953), .ZN(issueqPacket2_o[143]) );
  INVX0 U614 ( .INP(n956), .ZN(issueqPacket2_o[144]) );
  INVX0 U615 ( .INP(n1033), .ZN(issueqPacket1_o[37]) );
  INVX0 U616 ( .INP(n1036), .ZN(issueqPacket1_o[38]) );
  INVX0 U617 ( .INP(n1039), .ZN(issueqPacket1_o[39]) );
  INVX0 U618 ( .INP(n1042), .ZN(issueqPacket1_o[40]) );
  INVX0 U619 ( .INP(n1045), .ZN(issueqPacket1_o[41]) );
  INVX0 U620 ( .INP(n1048), .ZN(issueqPacket1_o[42]) );
  INVX0 U621 ( .INP(n1051), .ZN(issueqPacket1_o[43]) );
  INVX0 U622 ( .INP(n1054), .ZN(issueqPacket1_o[44]) );
  INVX0 U623 ( .INP(n1057), .ZN(issueqPacket1_o[45]) );
  INVX0 U624 ( .INP(n1060), .ZN(issueqPacket1_o[46]) );
  INVX0 U625 ( .INP(n1063), .ZN(issueqPacket1_o[47]) );
  INVX0 U626 ( .INP(n1066), .ZN(issueqPacket1_o[48]) );
  INVX0 U627 ( .INP(n1069), .ZN(issueqPacket1_o[49]) );
  INVX0 U628 ( .INP(n1072), .ZN(issueqPacket1_o[50]) );
  INVX0 U629 ( .INP(n1075), .ZN(issueqPacket1_o[51]) );
  INVX0 U630 ( .INP(n1078), .ZN(issueqPacket1_o[52]) );
  INVX0 U631 ( .INP(n1081), .ZN(issueqPacket1_o[53]) );
  INVX0 U632 ( .INP(n1084), .ZN(issueqPacket1_o[54]) );
  INVX0 U633 ( .INP(n1087), .ZN(issueqPacket1_o[55]) );
  INVX0 U634 ( .INP(n1090), .ZN(issueqPacket1_o[56]) );
  INVX0 U635 ( .INP(n1093), .ZN(issueqPacket1_o[57]) );
  INVX0 U636 ( .INP(n1096), .ZN(issueqPacket1_o[58]) );
  INVX0 U637 ( .INP(n1099), .ZN(issueqPacket1_o[59]) );
  INVX0 U638 ( .INP(n1102), .ZN(issueqPacket1_o[60]) );
  INVX0 U639 ( .INP(n1105), .ZN(issueqPacket1_o[61]) );
  INVX0 U640 ( .INP(n1108), .ZN(issueqPacket1_o[62]) );
  INVX0 U641 ( .INP(n1111), .ZN(issueqPacket1_o[63]) );
  INVX0 U642 ( .INP(n1114), .ZN(issueqPacket1_o[64]) );
  INVX0 U643 ( .INP(n1117), .ZN(issueqPacket1_o[65]) );
  INVX0 U644 ( .INP(n1120), .ZN(issueqPacket1_o[66]) );
  INVX0 U645 ( .INP(n1123), .ZN(issueqPacket1_o[67]) );
  INVX0 U646 ( .INP(n1126), .ZN(issueqPacket1_o[68]) );
  INVX0 U647 ( .INP(n1219), .ZN(issueqPacket1_o[114]) );
  INVX0 U648 ( .INP(n1222), .ZN(issueqPacket1_o[115]) );
  INVX0 U649 ( .INP(n1225), .ZN(issueqPacket1_o[116]) );
  INVX0 U650 ( .INP(n1228), .ZN(issueqPacket1_o[117]) );
  INVX0 U651 ( .INP(n1231), .ZN(issueqPacket1_o[118]) );
  INVX0 U652 ( .INP(n1234), .ZN(issueqPacket1_o[119]) );
  INVX0 U653 ( .INP(n1237), .ZN(issueqPacket1_o[120]) );
  INVX0 U654 ( .INP(n1240), .ZN(issueqPacket1_o[121]) );
  INVX0 U655 ( .INP(n1245), .ZN(issueqPacket1_o[123]) );
  INVX0 U656 ( .INP(n1248), .ZN(issueqPacket1_o[124]) );
  INVX0 U657 ( .INP(n1251), .ZN(issueqPacket1_o[125]) );
  INVX0 U658 ( .INP(n1254), .ZN(issueqPacket1_o[126]) );
  INVX0 U659 ( .INP(n1257), .ZN(issueqPacket1_o[127]) );
  INVX0 U660 ( .INP(n1260), .ZN(issueqPacket1_o[128]) );
  INVX0 U661 ( .INP(n1263), .ZN(issueqPacket1_o[129]) );
  INVX0 U662 ( .INP(n1280), .ZN(issueqPacket1_o[139]) );
  INVX0 U663 ( .INP(n1283), .ZN(issueqPacket1_o[140]) );
  INVX0 U664 ( .INP(n1286), .ZN(issueqPacket1_o[141]) );
  INVX0 U665 ( .INP(n1289), .ZN(issueqPacket1_o[142]) );
  INVX0 U666 ( .INP(n1292), .ZN(issueqPacket1_o[143]) );
  INVX0 U667 ( .INP(n1295), .ZN(issueqPacket1_o[144]) );
  INVX0 U668 ( .INP(n185), .ZN(issueqPacket0_o[37]) );
  INVX0 U669 ( .INP(n188), .ZN(issueqPacket0_o[38]) );
  INVX0 U670 ( .INP(n191), .ZN(issueqPacket0_o[39]) );
  INVX0 U671 ( .INP(n194), .ZN(issueqPacket0_o[40]) );
  INVX0 U672 ( .INP(n197), .ZN(issueqPacket0_o[41]) );
  INVX0 U673 ( .INP(n200), .ZN(issueqPacket0_o[42]) );
  INVX0 U674 ( .INP(n203), .ZN(issueqPacket0_o[43]) );
  INVX0 U675 ( .INP(n206), .ZN(issueqPacket0_o[44]) );
  INVX0 U676 ( .INP(n209), .ZN(issueqPacket0_o[45]) );
  INVX0 U677 ( .INP(n212), .ZN(issueqPacket0_o[46]) );
  INVX0 U678 ( .INP(n215), .ZN(issueqPacket0_o[47]) );
  INVX0 U679 ( .INP(n218), .ZN(issueqPacket0_o[48]) );
  INVX0 U680 ( .INP(n221), .ZN(issueqPacket0_o[49]) );
  INVX0 U681 ( .INP(n224), .ZN(issueqPacket0_o[50]) );
  INVX0 U682 ( .INP(n227), .ZN(issueqPacket0_o[51]) );
  INVX0 U683 ( .INP(n230), .ZN(issueqPacket0_o[52]) );
  INVX0 U684 ( .INP(n233), .ZN(issueqPacket0_o[53]) );
  INVX0 U685 ( .INP(n236), .ZN(issueqPacket0_o[54]) );
  INVX0 U686 ( .INP(n239), .ZN(issueqPacket0_o[55]) );
  INVX0 U687 ( .INP(n242), .ZN(issueqPacket0_o[56]) );
  INVX0 U688 ( .INP(n245), .ZN(issueqPacket0_o[57]) );
  INVX0 U689 ( .INP(n248), .ZN(issueqPacket0_o[58]) );
  INVX0 U690 ( .INP(n251), .ZN(issueqPacket0_o[59]) );
  INVX0 U691 ( .INP(n254), .ZN(issueqPacket0_o[60]) );
  INVX0 U692 ( .INP(n257), .ZN(issueqPacket0_o[61]) );
  INVX0 U693 ( .INP(n260), .ZN(issueqPacket0_o[62]) );
  INVX0 U694 ( .INP(n263), .ZN(issueqPacket0_o[63]) );
  INVX0 U695 ( .INP(n266), .ZN(issueqPacket0_o[64]) );
  INVX0 U696 ( .INP(n269), .ZN(issueqPacket0_o[65]) );
  INVX0 U697 ( .INP(n272), .ZN(issueqPacket0_o[66]) );
  INVX0 U698 ( .INP(n275), .ZN(issueqPacket0_o[67]) );
  INVX0 U699 ( .INP(n278), .ZN(issueqPacket0_o[68]) );
  INVX0 U700 ( .INP(n122), .ZN(issueqPacket0_o[114]) );
  INVX0 U701 ( .INP(n146), .ZN(issueqPacket0_o[115]) );
  INVX0 U702 ( .INP(n149), .ZN(issueqPacket0_o[116]) );
  INVX0 U703 ( .INP(n152), .ZN(issueqPacket0_o[117]) );
  INVX0 U704 ( .INP(n155), .ZN(issueqPacket0_o[118]) );
  INVX0 U705 ( .INP(n158), .ZN(issueqPacket0_o[119]) );
  INVX0 U706 ( .INP(n161), .ZN(issueqPacket0_o[120]) );
  INVX0 U707 ( .INP(n164), .ZN(issueqPacket0_o[121]) );
  INVX0 U708 ( .INP(n125), .ZN(issueqPacket0_o[123]) );
  INVX0 U709 ( .INP(n128), .ZN(issueqPacket0_o[124]) );
  INVX0 U710 ( .INP(n131), .ZN(issueqPacket0_o[125]) );
  INVX0 U711 ( .INP(n134), .ZN(issueqPacket0_o[126]) );
  INVX0 U712 ( .INP(n137), .ZN(issueqPacket0_o[127]) );
  INVX0 U713 ( .INP(n140), .ZN(issueqPacket0_o[128]) );
  INVX0 U714 ( .INP(n143), .ZN(issueqPacket0_o[129]) );
  INVX0 U715 ( .INP(n167), .ZN(issueqPacket0_o[139]) );
  INVX0 U716 ( .INP(n170), .ZN(issueqPacket0_o[140]) );
  INVX0 U717 ( .INP(n173), .ZN(issueqPacket0_o[141]) );
  INVX0 U718 ( .INP(n176), .ZN(issueqPacket0_o[142]) );
  INVX0 U719 ( .INP(n179), .ZN(issueqPacket0_o[143]) );
  INVX0 U720 ( .INP(n182), .ZN(issueqPacket0_o[144]) );
  INVX0 U721 ( .INP(ctrlVerifiedSMTid_i[1]), .ZN(n1478) );
  INVX0 U722 ( .INP(ctrlVerifiedSMTid_i[0]), .ZN(n1479) );
  INVX0 U723 ( .INP(n289), .ZN(issueqPacket3_o[0]) );
  INVX0 U724 ( .INP(renamedPacket3_i[0]), .ZN(n289) );
  INVX0 U725 ( .INP(n291), .ZN(issueqPacket3_o[1]) );
  INVX0 U726 ( .INP(renamedPacket3_i[1]), .ZN(n291) );
  INVX0 U727 ( .INP(n293), .ZN(issueqPacket3_o[2]) );
  INVX0 U728 ( .INP(renamedPacket3_i[2]), .ZN(n293) );
  INVX0 U729 ( .INP(n295), .ZN(issueqPacket3_o[3]) );
  INVX0 U730 ( .INP(renamedPacket3_i[3]), .ZN(n295) );
  INVX0 U731 ( .INP(n297), .ZN(issueqPacket3_o[4]) );
  INVX0 U732 ( .INP(renamedPacket3_i[4]), .ZN(n297) );
  INVX0 U733 ( .INP(n299), .ZN(issueqPacket3_o[5]) );
  INVX0 U734 ( .INP(renamedPacket3_i[5]), .ZN(n299) );
  INVX0 U735 ( .INP(n301), .ZN(issueqPacket3_o[6]) );
  INVX0 U736 ( .INP(renamedPacket3_i[6]), .ZN(n301) );
  INVX0 U737 ( .INP(n303), .ZN(issueqPacket3_o[7]) );
  INVX0 U738 ( .INP(renamedPacket3_i[7]), .ZN(n303) );
  INVX0 U739 ( .INP(n305), .ZN(issueqPacket3_o[8]) );
  INVX0 U740 ( .INP(renamedPacket3_i[8]), .ZN(n305) );
  INVX0 U741 ( .INP(n307), .ZN(issueqPacket3_o[9]) );
  INVX0 U742 ( .INP(renamedPacket3_i[9]), .ZN(n307) );
  INVX0 U743 ( .INP(n309), .ZN(issueqPacket3_o[10]) );
  INVX0 U744 ( .INP(renamedPacket3_i[10]), .ZN(n309) );
  INVX0 U745 ( .INP(n311), .ZN(issueqPacket3_o[11]) );
  INVX0 U746 ( .INP(renamedPacket3_i[11]), .ZN(n311) );
  INVX0 U747 ( .INP(n313), .ZN(issueqPacket3_o[12]) );
  INVX0 U748 ( .INP(renamedPacket3_i[12]), .ZN(n313) );
  INVX0 U749 ( .INP(n315), .ZN(issueqPacket3_o[13]) );
  INVX0 U750 ( .INP(renamedPacket3_i[13]), .ZN(n315) );
  INVX0 U751 ( .INP(n317), .ZN(issueqPacket3_o[14]) );
  INVX0 U752 ( .INP(renamedPacket3_i[14]), .ZN(n317) );
  INVX0 U753 ( .INP(n319), .ZN(issueqPacket3_o[15]) );
  INVX0 U754 ( .INP(renamedPacket3_i[15]), .ZN(n319) );
  INVX0 U755 ( .INP(n321), .ZN(issueqPacket3_o[16]) );
  INVX0 U756 ( .INP(renamedPacket3_i[16]), .ZN(n321) );
  INVX0 U757 ( .INP(n323), .ZN(issueqPacket3_o[17]) );
  INVX0 U758 ( .INP(renamedPacket3_i[17]), .ZN(n323) );
  INVX0 U759 ( .INP(n325), .ZN(issueqPacket3_o[18]) );
  INVX0 U760 ( .INP(renamedPacket3_i[18]), .ZN(n325) );
  INVX0 U761 ( .INP(n327), .ZN(issueqPacket3_o[19]) );
  INVX0 U762 ( .INP(renamedPacket3_i[19]), .ZN(n327) );
  INVX0 U763 ( .INP(n329), .ZN(issueqPacket3_o[20]) );
  INVX0 U764 ( .INP(renamedPacket3_i[20]), .ZN(n329) );
  INVX0 U765 ( .INP(n331), .ZN(issueqPacket3_o[21]) );
  INVX0 U766 ( .INP(renamedPacket3_i[21]), .ZN(n331) );
  INVX0 U767 ( .INP(n333), .ZN(issueqPacket3_o[22]) );
  INVX0 U768 ( .INP(renamedPacket3_i[22]), .ZN(n333) );
  INVX0 U769 ( .INP(n335), .ZN(issueqPacket3_o[23]) );
  INVX0 U770 ( .INP(renamedPacket3_i[23]), .ZN(n335) );
  INVX0 U771 ( .INP(n337), .ZN(issueqPacket3_o[24]) );
  INVX0 U772 ( .INP(renamedPacket3_i[24]), .ZN(n337) );
  INVX0 U773 ( .INP(n339), .ZN(issueqPacket3_o[25]) );
  INVX0 U774 ( .INP(renamedPacket3_i[25]), .ZN(n339) );
  INVX0 U775 ( .INP(n341), .ZN(issueqPacket3_o[26]) );
  INVX0 U776 ( .INP(renamedPacket3_i[26]), .ZN(n341) );
  INVX0 U777 ( .INP(n343), .ZN(issueqPacket3_o[27]) );
  INVX0 U778 ( .INP(renamedPacket3_i[27]), .ZN(n343) );
  INVX0 U779 ( .INP(n345), .ZN(issueqPacket3_o[28]) );
  INVX0 U780 ( .INP(renamedPacket3_i[28]), .ZN(n345) );
  INVX0 U781 ( .INP(n347), .ZN(issueqPacket3_o[29]) );
  INVX0 U782 ( .INP(renamedPacket3_i[29]), .ZN(n347) );
  INVX0 U783 ( .INP(n349), .ZN(issueqPacket3_o[30]) );
  INVX0 U784 ( .INP(renamedPacket3_i[30]), .ZN(n349) );
  INVX0 U785 ( .INP(n351), .ZN(issueqPacket3_o[31]) );
  INVX0 U786 ( .INP(renamedPacket3_i[31]), .ZN(n351) );
  INVX0 U787 ( .INP(n353), .ZN(issueqPacket3_o[32]) );
  INVX0 U788 ( .INP(renamedPacket3_i[32]), .ZN(n353) );
  INVX0 U789 ( .INP(n355), .ZN(issueqPacket3_o[33]) );
  INVX0 U790 ( .INP(renamedPacket3_i[33]), .ZN(n355) );
  INVX0 U791 ( .INP(n357), .ZN(issueqPacket3_o[34]) );
  INVX0 U792 ( .INP(renamedPacket3_i[34]), .ZN(n357) );
  INVX0 U793 ( .INP(n359), .ZN(issueqPacket3_o[35]) );
  INVX0 U794 ( .INP(renamedPacket3_i[35]), .ZN(n359) );
  INVX0 U795 ( .INP(n361), .ZN(issueqPacket3_o[36]) );
  INVX0 U796 ( .INP(renamedPacket3_i[36]), .ZN(n361) );
  INVX0 U797 ( .INP(n461), .ZN(issueqPacket3_o[70]) );
  INVX0 U798 ( .INP(renamedPacket3_i[70]), .ZN(n461) );
  INVX0 U799 ( .INP(n463), .ZN(issueqPacket3_o[71]) );
  INVX0 U800 ( .INP(renamedPacket3_i[71]), .ZN(n463) );
  INVX0 U801 ( .INP(n465), .ZN(issueqPacket3_o[72]) );
  INVX0 U802 ( .INP(renamedPacket3_i[72]), .ZN(n465) );
  INVX0 U803 ( .INP(n467), .ZN(issueqPacket3_o[73]) );
  INVX0 U804 ( .INP(renamedPacket3_i[73]), .ZN(n467) );
  INVX0 U805 ( .INP(n469), .ZN(issueqPacket3_o[74]) );
  INVX0 U806 ( .INP(renamedPacket3_i[74]), .ZN(n469) );
  INVX0 U807 ( .INP(n471), .ZN(issueqPacket3_o[75]) );
  INVX0 U808 ( .INP(renamedPacket3_i[75]), .ZN(n471) );
  INVX0 U809 ( .INP(n473), .ZN(issueqPacket3_o[76]) );
  INVX0 U810 ( .INP(renamedPacket3_i[76]), .ZN(n473) );
  INVX0 U811 ( .INP(n475), .ZN(issueqPacket3_o[77]) );
  INVX0 U812 ( .INP(renamedPacket3_i[77]), .ZN(n475) );
  INVX0 U813 ( .INP(n477), .ZN(issueqPacket3_o[78]) );
  INVX0 U814 ( .INP(renamedPacket3_i[78]), .ZN(n477) );
  INVX0 U815 ( .INP(n479), .ZN(issueqPacket3_o[79]) );
  INVX0 U816 ( .INP(renamedPacket3_i[79]), .ZN(n479) );
  INVX0 U817 ( .INP(n481), .ZN(issueqPacket3_o[80]) );
  INVX0 U818 ( .INP(renamedPacket3_i[80]), .ZN(n481) );
  INVX0 U819 ( .INP(n483), .ZN(issueqPacket3_o[81]) );
  INVX0 U820 ( .INP(renamedPacket3_i[81]), .ZN(n483) );
  INVX0 U821 ( .INP(n485), .ZN(issueqPacket3_o[82]) );
  INVX0 U822 ( .INP(renamedPacket3_i[82]), .ZN(n485) );
  INVX0 U823 ( .INP(n487), .ZN(issueqPacket3_o[83]) );
  INVX0 U824 ( .INP(renamedPacket3_i[83]), .ZN(n487) );
  INVX0 U825 ( .INP(n489), .ZN(issueqPacket3_o[84]) );
  INVX0 U826 ( .INP(renamedPacket3_i[84]), .ZN(n489) );
  INVX0 U827 ( .INP(n491), .ZN(issueqPacket3_o[85]) );
  INVX0 U828 ( .INP(renamedPacket3_i[85]), .ZN(n491) );
  INVX0 U829 ( .INP(n493), .ZN(issueqPacket3_o[86]) );
  INVX0 U830 ( .INP(renamedPacket3_i[86]), .ZN(n493) );
  INVX0 U831 ( .INP(n495), .ZN(issueqPacket3_o[87]) );
  INVX0 U832 ( .INP(renamedPacket3_i[87]), .ZN(n495) );
  INVX0 U833 ( .INP(n497), .ZN(issueqPacket3_o[88]) );
  INVX0 U834 ( .INP(renamedPacket3_i[88]), .ZN(n497) );
  INVX0 U835 ( .INP(n499), .ZN(issueqPacket3_o[89]) );
  INVX0 U836 ( .INP(renamedPacket3_i[89]), .ZN(n499) );
  INVX0 U837 ( .INP(n501), .ZN(issueqPacket3_o[90]) );
  INVX0 U838 ( .INP(renamedPacket3_i[90]), .ZN(n501) );
  INVX0 U839 ( .INP(n503), .ZN(issueqPacket3_o[91]) );
  INVX0 U840 ( .INP(renamedPacket3_i[91]), .ZN(n503) );
  INVX0 U841 ( .INP(n505), .ZN(issueqPacket3_o[92]) );
  INVX0 U842 ( .INP(renamedPacket3_i[92]), .ZN(n505) );
  INVX0 U843 ( .INP(n507), .ZN(issueqPacket3_o[93]) );
  INVX0 U844 ( .INP(renamedPacket3_i[93]), .ZN(n507) );
  INVX0 U845 ( .INP(n509), .ZN(issueqPacket3_o[94]) );
  INVX0 U846 ( .INP(renamedPacket3_i[94]), .ZN(n509) );
  INVX0 U847 ( .INP(n511), .ZN(issueqPacket3_o[95]) );
  INVX0 U848 ( .INP(renamedPacket3_i[95]), .ZN(n511) );
  INVX0 U849 ( .INP(n513), .ZN(issueqPacket3_o[96]) );
  INVX0 U850 ( .INP(renamedPacket3_i[96]), .ZN(n513) );
  INVX0 U851 ( .INP(n515), .ZN(issueqPacket3_o[97]) );
  INVX0 U852 ( .INP(renamedPacket3_i[97]), .ZN(n515) );
  INVX0 U853 ( .INP(n517), .ZN(issueqPacket3_o[98]) );
  INVX0 U854 ( .INP(renamedPacket3_i[98]), .ZN(n517) );
  INVX0 U855 ( .INP(n519), .ZN(issueqPacket3_o[99]) );
  INVX0 U856 ( .INP(renamedPacket3_i[99]), .ZN(n519) );
  INVX0 U857 ( .INP(n521), .ZN(issueqPacket3_o[100]) );
  INVX0 U858 ( .INP(renamedPacket3_i[100]), .ZN(n521) );
  INVX0 U859 ( .INP(n523), .ZN(issueqPacket3_o[101]) );
  INVX0 U860 ( .INP(renamedPacket3_i[101]), .ZN(n523) );
  INVX0 U861 ( .INP(n525), .ZN(issueqPacket3_o[102]) );
  INVX0 U862 ( .INP(renamedPacket3_i[102]), .ZN(n525) );
  INVX0 U863 ( .INP(n527), .ZN(issueqPacket3_o[103]) );
  INVX0 U864 ( .INP(renamedPacket3_i[103]), .ZN(n527) );
  INVX0 U865 ( .INP(n529), .ZN(issueqPacket3_o[104]) );
  INVX0 U866 ( .INP(renamedPacket3_i[104]), .ZN(n529) );
  INVX0 U867 ( .INP(n531), .ZN(issueqPacket3_o[105]) );
  INVX0 U868 ( .INP(renamedPacket3_i[105]), .ZN(n531) );
  INVX0 U869 ( .INP(n533), .ZN(issueqPacket3_o[106]) );
  INVX0 U870 ( .INP(renamedPacket3_i[106]), .ZN(n533) );
  INVX0 U871 ( .INP(n535), .ZN(issueqPacket3_o[107]) );
  INVX0 U872 ( .INP(renamedPacket3_i[107]), .ZN(n535) );
  INVX0 U873 ( .INP(n537), .ZN(issueqPacket3_o[108]) );
  INVX0 U874 ( .INP(renamedPacket3_i[108]), .ZN(n537) );
  INVX0 U875 ( .INP(n539), .ZN(issueqPacket3_o[109]) );
  INVX0 U876 ( .INP(renamedPacket3_i[109]), .ZN(n539) );
  INVX0 U877 ( .INP(n541), .ZN(issueqPacket3_o[110]) );
  INVX0 U878 ( .INP(renamedPacket3_i[110]), .ZN(n541) );
  INVX0 U879 ( .INP(n543), .ZN(issueqPacket3_o[111]) );
  INVX0 U880 ( .INP(renamedPacket3_i[111]), .ZN(n543) );
  INVX0 U881 ( .INP(n545), .ZN(issueqPacket3_o[112]) );
  INVX0 U882 ( .INP(renamedPacket3_i[112]), .ZN(n545) );
  INVX0 U883 ( .INP(n547), .ZN(issueqPacket3_o[113]) );
  INVX0 U884 ( .INP(renamedPacket3_i[113]), .ZN(n547) );
  INVX0 U885 ( .INP(n573), .ZN(issueqPacket3_o[122]) );
  INVX0 U886 ( .INP(renamedPacket3_i[122]), .ZN(n573) );
  INVX0 U887 ( .INP(n596), .ZN(issueqPacket3_o[130]) );
  INVX0 U888 ( .INP(renamedPacket3_i[130]), .ZN(n596) );
  INVX0 U889 ( .INP(n598), .ZN(issueqPacket3_o[131]) );
  INVX0 U890 ( .INP(renamedPacket3_i[131]), .ZN(n598) );
  INVX0 U891 ( .INP(n600), .ZN(issueqPacket3_o[138]) );
  INVX0 U892 ( .INP(issueqPacket3_o_138), .ZN(n600) );
  INVX0 U893 ( .INP(n620), .ZN(issueqPacket2_o[0]) );
  INVX0 U894 ( .INP(renamedPacket2_i[0]), .ZN(n620) );
  INVX0 U895 ( .INP(n622), .ZN(issueqPacket2_o[1]) );
  INVX0 U896 ( .INP(renamedPacket2_i[1]), .ZN(n622) );
  INVX0 U897 ( .INP(n624), .ZN(issueqPacket2_o[2]) );
  INVX0 U898 ( .INP(renamedPacket2_i[2]), .ZN(n624) );
  INVX0 U899 ( .INP(n626), .ZN(issueqPacket2_o[3]) );
  INVX0 U900 ( .INP(renamedPacket2_i[3]), .ZN(n626) );
  INVX0 U901 ( .INP(n628), .ZN(issueqPacket2_o[4]) );
  INVX0 U902 ( .INP(renamedPacket2_i[4]), .ZN(n628) );
  INVX0 U903 ( .INP(n630), .ZN(issueqPacket2_o[5]) );
  INVX0 U904 ( .INP(renamedPacket2_i[5]), .ZN(n630) );
  INVX0 U905 ( .INP(n632), .ZN(issueqPacket2_o[6]) );
  INVX0 U906 ( .INP(renamedPacket2_i[6]), .ZN(n632) );
  INVX0 U907 ( .INP(n634), .ZN(issueqPacket2_o[7]) );
  INVX0 U908 ( .INP(renamedPacket2_i[7]), .ZN(n634) );
  INVX0 U909 ( .INP(n636), .ZN(issueqPacket2_o[8]) );
  INVX0 U910 ( .INP(renamedPacket2_i[8]), .ZN(n636) );
  INVX0 U911 ( .INP(n638), .ZN(issueqPacket2_o[9]) );
  INVX0 U912 ( .INP(renamedPacket2_i[9]), .ZN(n638) );
  INVX0 U913 ( .INP(n640), .ZN(issueqPacket2_o[10]) );
  INVX0 U914 ( .INP(renamedPacket2_i[10]), .ZN(n640) );
  INVX0 U915 ( .INP(n642), .ZN(issueqPacket2_o[11]) );
  INVX0 U916 ( .INP(renamedPacket2_i[11]), .ZN(n642) );
  INVX0 U917 ( .INP(n644), .ZN(issueqPacket2_o[12]) );
  INVX0 U918 ( .INP(renamedPacket2_i[12]), .ZN(n644) );
  INVX0 U919 ( .INP(n646), .ZN(issueqPacket2_o[13]) );
  INVX0 U920 ( .INP(renamedPacket2_i[13]), .ZN(n646) );
  INVX0 U921 ( .INP(n648), .ZN(issueqPacket2_o[14]) );
  INVX0 U922 ( .INP(renamedPacket2_i[14]), .ZN(n648) );
  INVX0 U923 ( .INP(n650), .ZN(issueqPacket2_o[15]) );
  INVX0 U924 ( .INP(renamedPacket2_i[15]), .ZN(n650) );
  INVX0 U925 ( .INP(n652), .ZN(issueqPacket2_o[16]) );
  INVX0 U926 ( .INP(renamedPacket2_i[16]), .ZN(n652) );
  INVX0 U927 ( .INP(n654), .ZN(issueqPacket2_o[17]) );
  INVX0 U928 ( .INP(renamedPacket2_i[17]), .ZN(n654) );
  INVX0 U929 ( .INP(n656), .ZN(issueqPacket2_o[18]) );
  INVX0 U930 ( .INP(renamedPacket2_i[18]), .ZN(n656) );
  INVX0 U931 ( .INP(n658), .ZN(issueqPacket2_o[19]) );
  INVX0 U932 ( .INP(renamedPacket2_i[19]), .ZN(n658) );
  INVX0 U933 ( .INP(n660), .ZN(issueqPacket2_o[20]) );
  INVX0 U934 ( .INP(renamedPacket2_i[20]), .ZN(n660) );
  INVX0 U935 ( .INP(n662), .ZN(issueqPacket2_o[21]) );
  INVX0 U936 ( .INP(renamedPacket2_i[21]), .ZN(n662) );
  INVX0 U937 ( .INP(n664), .ZN(issueqPacket2_o[22]) );
  INVX0 U938 ( .INP(renamedPacket2_i[22]), .ZN(n664) );
  INVX0 U939 ( .INP(n666), .ZN(issueqPacket2_o[23]) );
  INVX0 U940 ( .INP(renamedPacket2_i[23]), .ZN(n666) );
  INVX0 U941 ( .INP(n668), .ZN(issueqPacket2_o[24]) );
  INVX0 U942 ( .INP(renamedPacket2_i[24]), .ZN(n668) );
  INVX0 U943 ( .INP(n670), .ZN(issueqPacket2_o[25]) );
  INVX0 U944 ( .INP(renamedPacket2_i[25]), .ZN(n670) );
  INVX0 U945 ( .INP(n672), .ZN(issueqPacket2_o[26]) );
  INVX0 U946 ( .INP(renamedPacket2_i[26]), .ZN(n672) );
  INVX0 U947 ( .INP(n674), .ZN(issueqPacket2_o[27]) );
  INVX0 U948 ( .INP(renamedPacket2_i[27]), .ZN(n674) );
  INVX0 U949 ( .INP(n676), .ZN(issueqPacket2_o[28]) );
  INVX0 U950 ( .INP(renamedPacket2_i[28]), .ZN(n676) );
  INVX0 U951 ( .INP(n678), .ZN(issueqPacket2_o[29]) );
  INVX0 U952 ( .INP(renamedPacket2_i[29]), .ZN(n678) );
  INVX0 U953 ( .INP(n680), .ZN(issueqPacket2_o[30]) );
  INVX0 U954 ( .INP(renamedPacket2_i[30]), .ZN(n680) );
  INVX0 U955 ( .INP(n682), .ZN(issueqPacket2_o[31]) );
  INVX0 U956 ( .INP(renamedPacket2_i[31]), .ZN(n682) );
  INVX0 U957 ( .INP(n684), .ZN(issueqPacket2_o[32]) );
  INVX0 U958 ( .INP(renamedPacket2_i[32]), .ZN(n684) );
  INVX0 U959 ( .INP(n686), .ZN(issueqPacket2_o[33]) );
  INVX0 U960 ( .INP(renamedPacket2_i[33]), .ZN(n686) );
  INVX0 U961 ( .INP(n688), .ZN(issueqPacket2_o[34]) );
  INVX0 U962 ( .INP(renamedPacket2_i[34]), .ZN(n688) );
  INVX0 U963 ( .INP(n690), .ZN(issueqPacket2_o[35]) );
  INVX0 U964 ( .INP(renamedPacket2_i[35]), .ZN(n690) );
  INVX0 U965 ( .INP(n692), .ZN(issueqPacket2_o[36]) );
  INVX0 U966 ( .INP(renamedPacket2_i[36]), .ZN(n692) );
  INVX0 U967 ( .INP(n790), .ZN(issueqPacket2_o[69]) );
  INVX0 U968 ( .INP(renamedPacket2_i[69]), .ZN(n790) );
  INVX0 U969 ( .INP(n792), .ZN(issueqPacket2_o[70]) );
  INVX0 U970 ( .INP(renamedPacket2_i[70]), .ZN(n792) );
  INVX0 U971 ( .INP(n794), .ZN(issueqPacket2_o[71]) );
  INVX0 U972 ( .INP(renamedPacket2_i[71]), .ZN(n794) );
  INVX0 U973 ( .INP(n796), .ZN(issueqPacket2_o[72]) );
  INVX0 U974 ( .INP(renamedPacket2_i[72]), .ZN(n796) );
  INVX0 U975 ( .INP(n798), .ZN(issueqPacket2_o[73]) );
  INVX0 U976 ( .INP(renamedPacket2_i[73]), .ZN(n798) );
  INVX0 U977 ( .INP(n800), .ZN(issueqPacket2_o[74]) );
  INVX0 U978 ( .INP(renamedPacket2_i[74]), .ZN(n800) );
  INVX0 U979 ( .INP(n802), .ZN(issueqPacket2_o[75]) );
  INVX0 U980 ( .INP(renamedPacket2_i[75]), .ZN(n802) );
  INVX0 U981 ( .INP(n804), .ZN(issueqPacket2_o[76]) );
  INVX0 U982 ( .INP(renamedPacket2_i[76]), .ZN(n804) );
  INVX0 U983 ( .INP(n806), .ZN(issueqPacket2_o[77]) );
  INVX0 U984 ( .INP(renamedPacket2_i[77]), .ZN(n806) );
  INVX0 U985 ( .INP(n808), .ZN(issueqPacket2_o[78]) );
  INVX0 U986 ( .INP(renamedPacket2_i[78]), .ZN(n808) );
  INVX0 U987 ( .INP(n810), .ZN(issueqPacket2_o[79]) );
  INVX0 U988 ( .INP(renamedPacket2_i[79]), .ZN(n810) );
  INVX0 U989 ( .INP(n812), .ZN(issueqPacket2_o[80]) );
  INVX0 U990 ( .INP(renamedPacket2_i[80]), .ZN(n812) );
  INVX0 U991 ( .INP(n814), .ZN(issueqPacket2_o[81]) );
  INVX0 U992 ( .INP(renamedPacket2_i[81]), .ZN(n814) );
  INVX0 U993 ( .INP(n816), .ZN(issueqPacket2_o[82]) );
  INVX0 U994 ( .INP(renamedPacket2_i[82]), .ZN(n816) );
  INVX0 U995 ( .INP(n818), .ZN(issueqPacket2_o[83]) );
  INVX0 U996 ( .INP(renamedPacket2_i[83]), .ZN(n818) );
  INVX0 U997 ( .INP(n820), .ZN(issueqPacket2_o[84]) );
  INVX0 U998 ( .INP(renamedPacket2_i[84]), .ZN(n820) );
  INVX0 U999 ( .INP(n822), .ZN(issueqPacket2_o[85]) );
  INVX0 U1000 ( .INP(renamedPacket2_i[85]), .ZN(n822) );
  INVX0 U1001 ( .INP(n824), .ZN(issueqPacket2_o[86]) );
  INVX0 U1002 ( .INP(renamedPacket2_i[86]), .ZN(n824) );
  INVX0 U1003 ( .INP(n826), .ZN(issueqPacket2_o[87]) );
  INVX0 U1004 ( .INP(renamedPacket2_i[87]), .ZN(n826) );
  INVX0 U1005 ( .INP(n828), .ZN(issueqPacket2_o[88]) );
  INVX0 U1006 ( .INP(renamedPacket2_i[88]), .ZN(n828) );
  INVX0 U1007 ( .INP(n830), .ZN(issueqPacket2_o[89]) );
  INVX0 U1008 ( .INP(renamedPacket2_i[89]), .ZN(n830) );
  INVX0 U1009 ( .INP(n832), .ZN(issueqPacket2_o[90]) );
  INVX0 U1010 ( .INP(renamedPacket2_i[90]), .ZN(n832) );
  INVX0 U1011 ( .INP(n834), .ZN(issueqPacket2_o[91]) );
  INVX0 U1012 ( .INP(renamedPacket2_i[91]), .ZN(n834) );
  INVX0 U1013 ( .INP(n836), .ZN(issueqPacket2_o[92]) );
  INVX0 U1014 ( .INP(renamedPacket2_i[92]), .ZN(n836) );
  INVX0 U1015 ( .INP(n838), .ZN(issueqPacket2_o[93]) );
  INVX0 U1016 ( .INP(renamedPacket2_i[93]), .ZN(n838) );
  INVX0 U1017 ( .INP(n840), .ZN(issueqPacket2_o[94]) );
  INVX0 U1018 ( .INP(renamedPacket2_i[94]), .ZN(n840) );
  INVX0 U1019 ( .INP(n842), .ZN(issueqPacket2_o[95]) );
  INVX0 U1020 ( .INP(renamedPacket2_i[95]), .ZN(n842) );
  INVX0 U1021 ( .INP(n844), .ZN(issueqPacket2_o[96]) );
  INVX0 U1022 ( .INP(renamedPacket2_i[96]), .ZN(n844) );
  INVX0 U1023 ( .INP(n846), .ZN(issueqPacket2_o[97]) );
  INVX0 U1024 ( .INP(renamedPacket2_i[97]), .ZN(n846) );
  INVX0 U1025 ( .INP(n848), .ZN(issueqPacket2_o[98]) );
  INVX0 U1026 ( .INP(renamedPacket2_i[98]), .ZN(n848) );
  INVX0 U1027 ( .INP(n850), .ZN(issueqPacket2_o[99]) );
  INVX0 U1028 ( .INP(renamedPacket2_i[99]), .ZN(n850) );
  INVX0 U1029 ( .INP(n852), .ZN(issueqPacket2_o[100]) );
  INVX0 U1030 ( .INP(renamedPacket2_i[100]), .ZN(n852) );
  INVX0 U1031 ( .INP(n854), .ZN(issueqPacket2_o[101]) );
  INVX0 U1032 ( .INP(renamedPacket2_i[101]), .ZN(n854) );
  INVX0 U1033 ( .INP(n856), .ZN(issueqPacket2_o[102]) );
  INVX0 U1034 ( .INP(renamedPacket2_i[102]), .ZN(n856) );
  INVX0 U1035 ( .INP(n858), .ZN(issueqPacket2_o[103]) );
  INVX0 U1036 ( .INP(renamedPacket2_i[103]), .ZN(n858) );
  INVX0 U1037 ( .INP(n860), .ZN(issueqPacket2_o[104]) );
  INVX0 U1038 ( .INP(renamedPacket2_i[104]), .ZN(n860) );
  INVX0 U1039 ( .INP(n862), .ZN(issueqPacket2_o[105]) );
  INVX0 U1040 ( .INP(renamedPacket2_i[105]), .ZN(n862) );
  INVX0 U1041 ( .INP(n864), .ZN(issueqPacket2_o[106]) );
  INVX0 U1042 ( .INP(renamedPacket2_i[106]), .ZN(n864) );
  INVX0 U1043 ( .INP(n866), .ZN(issueqPacket2_o[107]) );
  INVX0 U1044 ( .INP(renamedPacket2_i[107]), .ZN(n866) );
  INVX0 U1045 ( .INP(n868), .ZN(issueqPacket2_o[108]) );
  INVX0 U1046 ( .INP(renamedPacket2_i[108]), .ZN(n868) );
  INVX0 U1047 ( .INP(n870), .ZN(issueqPacket2_o[109]) );
  INVX0 U1048 ( .INP(renamedPacket2_i[109]), .ZN(n870) );
  INVX0 U1049 ( .INP(n872), .ZN(issueqPacket2_o[110]) );
  INVX0 U1050 ( .INP(renamedPacket2_i[110]), .ZN(n872) );
  INVX0 U1051 ( .INP(n874), .ZN(issueqPacket2_o[111]) );
  INVX0 U1052 ( .INP(renamedPacket2_i[111]), .ZN(n874) );
  INVX0 U1053 ( .INP(n876), .ZN(issueqPacket2_o[112]) );
  INVX0 U1054 ( .INP(renamedPacket2_i[112]), .ZN(n876) );
  INVX0 U1055 ( .INP(n878), .ZN(issueqPacket2_o[113]) );
  INVX0 U1056 ( .INP(renamedPacket2_i[113]), .ZN(n878) );
  INVX0 U1057 ( .INP(n904), .ZN(issueqPacket2_o[122]) );
  INVX0 U1058 ( .INP(renamedPacket2_i[122]), .ZN(n904) );
  INVX0 U1059 ( .INP(n927), .ZN(issueqPacket2_o[130]) );
  INVX0 U1060 ( .INP(renamedPacket2_i[130]), .ZN(n927) );
  INVX0 U1061 ( .INP(n929), .ZN(issueqPacket2_o[131]) );
  INVX0 U1062 ( .INP(renamedPacket2_i[131]), .ZN(n929) );
  INVX0 U1063 ( .INP(n939), .ZN(issueqPacket2_o[138]) );
  INVX0 U1064 ( .INP(issueqPacket2_o_138), .ZN(n939) );
  INVX0 U1065 ( .INP(n959), .ZN(issueqPacket1_o[0]) );
  INVX0 U1066 ( .INP(renamedPacket1_i[0]), .ZN(n959) );
  INVX0 U1067 ( .INP(n961), .ZN(issueqPacket1_o[1]) );
  INVX0 U1068 ( .INP(renamedPacket1_i[1]), .ZN(n961) );
  INVX0 U1069 ( .INP(n963), .ZN(issueqPacket1_o[2]) );
  INVX0 U1070 ( .INP(renamedPacket1_i[2]), .ZN(n963) );
  INVX0 U1071 ( .INP(n965), .ZN(issueqPacket1_o[3]) );
  INVX0 U1072 ( .INP(renamedPacket1_i[3]), .ZN(n965) );
  INVX0 U1073 ( .INP(n967), .ZN(issueqPacket1_o[4]) );
  INVX0 U1074 ( .INP(renamedPacket1_i[4]), .ZN(n967) );
  INVX0 U1075 ( .INP(n969), .ZN(issueqPacket1_o[5]) );
  INVX0 U1076 ( .INP(renamedPacket1_i[5]), .ZN(n969) );
  INVX0 U1077 ( .INP(n971), .ZN(issueqPacket1_o[6]) );
  INVX0 U1078 ( .INP(renamedPacket1_i[6]), .ZN(n971) );
  INVX0 U1079 ( .INP(n973), .ZN(issueqPacket1_o[7]) );
  INVX0 U1080 ( .INP(renamedPacket1_i[7]), .ZN(n973) );
  INVX0 U1081 ( .INP(n975), .ZN(issueqPacket1_o[8]) );
  INVX0 U1082 ( .INP(renamedPacket1_i[8]), .ZN(n975) );
  INVX0 U1083 ( .INP(n977), .ZN(issueqPacket1_o[9]) );
  INVX0 U1084 ( .INP(renamedPacket1_i[9]), .ZN(n977) );
  INVX0 U1085 ( .INP(n979), .ZN(issueqPacket1_o[10]) );
  INVX0 U1086 ( .INP(renamedPacket1_i[10]), .ZN(n979) );
  INVX0 U1087 ( .INP(n981), .ZN(issueqPacket1_o[11]) );
  INVX0 U1088 ( .INP(renamedPacket1_i[11]), .ZN(n981) );
  INVX0 U1089 ( .INP(n983), .ZN(issueqPacket1_o[12]) );
  INVX0 U1090 ( .INP(renamedPacket1_i[12]), .ZN(n983) );
  INVX0 U1091 ( .INP(n985), .ZN(issueqPacket1_o[13]) );
  INVX0 U1092 ( .INP(renamedPacket1_i[13]), .ZN(n985) );
  INVX0 U1093 ( .INP(n987), .ZN(issueqPacket1_o[14]) );
  INVX0 U1094 ( .INP(renamedPacket1_i[14]), .ZN(n987) );
  INVX0 U1095 ( .INP(n989), .ZN(issueqPacket1_o[15]) );
  INVX0 U1096 ( .INP(renamedPacket1_i[15]), .ZN(n989) );
  INVX0 U1097 ( .INP(n991), .ZN(issueqPacket1_o[16]) );
  INVX0 U1098 ( .INP(renamedPacket1_i[16]), .ZN(n991) );
  INVX0 U1099 ( .INP(n993), .ZN(issueqPacket1_o[17]) );
  INVX0 U1100 ( .INP(renamedPacket1_i[17]), .ZN(n993) );
  INVX0 U1101 ( .INP(n995), .ZN(issueqPacket1_o[18]) );
  INVX0 U1102 ( .INP(renamedPacket1_i[18]), .ZN(n995) );
  INVX0 U1103 ( .INP(n997), .ZN(issueqPacket1_o[19]) );
  INVX0 U1104 ( .INP(renamedPacket1_i[19]), .ZN(n997) );
  INVX0 U1105 ( .INP(n999), .ZN(issueqPacket1_o[20]) );
  INVX0 U1106 ( .INP(renamedPacket1_i[20]), .ZN(n999) );
  INVX0 U1107 ( .INP(n1001), .ZN(issueqPacket1_o[21]) );
  INVX0 U1108 ( .INP(renamedPacket1_i[21]), .ZN(n1001) );
  INVX0 U1109 ( .INP(n1003), .ZN(issueqPacket1_o[22]) );
  INVX0 U1110 ( .INP(renamedPacket1_i[22]), .ZN(n1003) );
  INVX0 U1111 ( .INP(n1005), .ZN(issueqPacket1_o[23]) );
  INVX0 U1112 ( .INP(renamedPacket1_i[23]), .ZN(n1005) );
  INVX0 U1113 ( .INP(n1007), .ZN(issueqPacket1_o[24]) );
  INVX0 U1114 ( .INP(renamedPacket1_i[24]), .ZN(n1007) );
  INVX0 U1115 ( .INP(n1009), .ZN(issueqPacket1_o[25]) );
  INVX0 U1116 ( .INP(renamedPacket1_i[25]), .ZN(n1009) );
  INVX0 U1117 ( .INP(n1011), .ZN(issueqPacket1_o[26]) );
  INVX0 U1118 ( .INP(renamedPacket1_i[26]), .ZN(n1011) );
  INVX0 U1119 ( .INP(n1013), .ZN(issueqPacket1_o[27]) );
  INVX0 U1120 ( .INP(renamedPacket1_i[27]), .ZN(n1013) );
  INVX0 U1121 ( .INP(n1015), .ZN(issueqPacket1_o[28]) );
  INVX0 U1122 ( .INP(renamedPacket1_i[28]), .ZN(n1015) );
  INVX0 U1123 ( .INP(n1017), .ZN(issueqPacket1_o[29]) );
  INVX0 U1124 ( .INP(renamedPacket1_i[29]), .ZN(n1017) );
  INVX0 U1125 ( .INP(n1019), .ZN(issueqPacket1_o[30]) );
  INVX0 U1126 ( .INP(renamedPacket1_i[30]), .ZN(n1019) );
  INVX0 U1127 ( .INP(n1021), .ZN(issueqPacket1_o[31]) );
  INVX0 U1128 ( .INP(renamedPacket1_i[31]), .ZN(n1021) );
  INVX0 U1129 ( .INP(n1023), .ZN(issueqPacket1_o[32]) );
  INVX0 U1130 ( .INP(renamedPacket1_i[32]), .ZN(n1023) );
  INVX0 U1131 ( .INP(n1025), .ZN(issueqPacket1_o[33]) );
  INVX0 U1132 ( .INP(renamedPacket1_i[33]), .ZN(n1025) );
  INVX0 U1133 ( .INP(n1027), .ZN(issueqPacket1_o[34]) );
  INVX0 U1134 ( .INP(renamedPacket1_i[34]), .ZN(n1027) );
  INVX0 U1135 ( .INP(n1029), .ZN(issueqPacket1_o[35]) );
  INVX0 U1136 ( .INP(renamedPacket1_i[35]), .ZN(n1029) );
  INVX0 U1137 ( .INP(n1031), .ZN(issueqPacket1_o[36]) );
  INVX0 U1138 ( .INP(renamedPacket1_i[36]), .ZN(n1031) );
  INVX0 U1139 ( .INP(n1129), .ZN(issueqPacket1_o[69]) );
  INVX0 U1140 ( .INP(renamedPacket1_i[69]), .ZN(n1129) );
  INVX0 U1141 ( .INP(n1131), .ZN(issueqPacket1_o[70]) );
  INVX0 U1142 ( .INP(renamedPacket1_i[70]), .ZN(n1131) );
  INVX0 U1143 ( .INP(n1133), .ZN(issueqPacket1_o[71]) );
  INVX0 U1144 ( .INP(renamedPacket1_i[71]), .ZN(n1133) );
  INVX0 U1145 ( .INP(n1135), .ZN(issueqPacket1_o[72]) );
  INVX0 U1146 ( .INP(renamedPacket1_i[72]), .ZN(n1135) );
  INVX0 U1147 ( .INP(n1137), .ZN(issueqPacket1_o[73]) );
  INVX0 U1148 ( .INP(renamedPacket1_i[73]), .ZN(n1137) );
  INVX0 U1149 ( .INP(n1139), .ZN(issueqPacket1_o[74]) );
  INVX0 U1150 ( .INP(renamedPacket1_i[74]), .ZN(n1139) );
  INVX0 U1151 ( .INP(n1141), .ZN(issueqPacket1_o[75]) );
  INVX0 U1152 ( .INP(renamedPacket1_i[75]), .ZN(n1141) );
  INVX0 U1153 ( .INP(n1143), .ZN(issueqPacket1_o[76]) );
  INVX0 U1154 ( .INP(renamedPacket1_i[76]), .ZN(n1143) );
  INVX0 U1155 ( .INP(n1145), .ZN(issueqPacket1_o[77]) );
  INVX0 U1156 ( .INP(renamedPacket1_i[77]), .ZN(n1145) );
  INVX0 U1157 ( .INP(n1147), .ZN(issueqPacket1_o[78]) );
  INVX0 U1158 ( .INP(renamedPacket1_i[78]), .ZN(n1147) );
  INVX0 U1159 ( .INP(n1149), .ZN(issueqPacket1_o[79]) );
  INVX0 U1160 ( .INP(renamedPacket1_i[79]), .ZN(n1149) );
  INVX0 U1161 ( .INP(n1151), .ZN(issueqPacket1_o[80]) );
  INVX0 U1162 ( .INP(renamedPacket1_i[80]), .ZN(n1151) );
  INVX0 U1163 ( .INP(n1153), .ZN(issueqPacket1_o[81]) );
  INVX0 U1164 ( .INP(renamedPacket1_i[81]), .ZN(n1153) );
  INVX0 U1165 ( .INP(n1155), .ZN(issueqPacket1_o[82]) );
  INVX0 U1166 ( .INP(renamedPacket1_i[82]), .ZN(n1155) );
  INVX0 U1167 ( .INP(n1157), .ZN(issueqPacket1_o[83]) );
  INVX0 U1168 ( .INP(renamedPacket1_i[83]), .ZN(n1157) );
  INVX0 U1169 ( .INP(n1159), .ZN(issueqPacket1_o[84]) );
  INVX0 U1170 ( .INP(renamedPacket1_i[84]), .ZN(n1159) );
  INVX0 U1171 ( .INP(n1161), .ZN(issueqPacket1_o[85]) );
  INVX0 U1172 ( .INP(renamedPacket1_i[85]), .ZN(n1161) );
  INVX0 U1173 ( .INP(n1163), .ZN(issueqPacket1_o[86]) );
  INVX0 U1174 ( .INP(renamedPacket1_i[86]), .ZN(n1163) );
  INVX0 U1175 ( .INP(n1165), .ZN(issueqPacket1_o[87]) );
  INVX0 U1176 ( .INP(renamedPacket1_i[87]), .ZN(n1165) );
  INVX0 U1177 ( .INP(n1167), .ZN(issueqPacket1_o[88]) );
  INVX0 U1178 ( .INP(renamedPacket1_i[88]), .ZN(n1167) );
  INVX0 U1179 ( .INP(n1169), .ZN(issueqPacket1_o[89]) );
  INVX0 U1180 ( .INP(renamedPacket1_i[89]), .ZN(n1169) );
  INVX0 U1181 ( .INP(n1171), .ZN(issueqPacket1_o[90]) );
  INVX0 U1182 ( .INP(renamedPacket1_i[90]), .ZN(n1171) );
  INVX0 U1183 ( .INP(n1173), .ZN(issueqPacket1_o[91]) );
  INVX0 U1184 ( .INP(renamedPacket1_i[91]), .ZN(n1173) );
  INVX0 U1185 ( .INP(n1175), .ZN(issueqPacket1_o[92]) );
  INVX0 U1186 ( .INP(renamedPacket1_i[92]), .ZN(n1175) );
  INVX0 U1187 ( .INP(n1177), .ZN(issueqPacket1_o[93]) );
  INVX0 U1188 ( .INP(renamedPacket1_i[93]), .ZN(n1177) );
  INVX0 U1189 ( .INP(n1179), .ZN(issueqPacket1_o[94]) );
  INVX0 U1190 ( .INP(renamedPacket1_i[94]), .ZN(n1179) );
  INVX0 U1191 ( .INP(n1181), .ZN(issueqPacket1_o[95]) );
  INVX0 U1192 ( .INP(renamedPacket1_i[95]), .ZN(n1181) );
  INVX0 U1193 ( .INP(n1183), .ZN(issueqPacket1_o[96]) );
  INVX0 U1194 ( .INP(renamedPacket1_i[96]), .ZN(n1183) );
  INVX0 U1195 ( .INP(n1185), .ZN(issueqPacket1_o[97]) );
  INVX0 U1196 ( .INP(renamedPacket1_i[97]), .ZN(n1185) );
  INVX0 U1197 ( .INP(n1187), .ZN(issueqPacket1_o[98]) );
  INVX0 U1198 ( .INP(renamedPacket1_i[98]), .ZN(n1187) );
  INVX0 U1199 ( .INP(n1189), .ZN(issueqPacket1_o[99]) );
  INVX0 U1200 ( .INP(renamedPacket1_i[99]), .ZN(n1189) );
  INVX0 U1201 ( .INP(n1191), .ZN(issueqPacket1_o[100]) );
  INVX0 U1202 ( .INP(renamedPacket1_i[100]), .ZN(n1191) );
  INVX0 U1203 ( .INP(n1193), .ZN(issueqPacket1_o[101]) );
  INVX0 U1204 ( .INP(renamedPacket1_i[101]), .ZN(n1193) );
  INVX0 U1205 ( .INP(n1195), .ZN(issueqPacket1_o[102]) );
  INVX0 U1206 ( .INP(renamedPacket1_i[102]), .ZN(n1195) );
  INVX0 U1207 ( .INP(n1197), .ZN(issueqPacket1_o[103]) );
  INVX0 U1208 ( .INP(renamedPacket1_i[103]), .ZN(n1197) );
  INVX0 U1209 ( .INP(n1199), .ZN(issueqPacket1_o[104]) );
  INVX0 U1210 ( .INP(renamedPacket1_i[104]), .ZN(n1199) );
  INVX0 U1211 ( .INP(n1201), .ZN(issueqPacket1_o[105]) );
  INVX0 U1212 ( .INP(renamedPacket1_i[105]), .ZN(n1201) );
  INVX0 U1213 ( .INP(n1203), .ZN(issueqPacket1_o[106]) );
  INVX0 U1214 ( .INP(renamedPacket1_i[106]), .ZN(n1203) );
  INVX0 U1215 ( .INP(n1205), .ZN(issueqPacket1_o[107]) );
  INVX0 U1216 ( .INP(renamedPacket1_i[107]), .ZN(n1205) );
  INVX0 U1217 ( .INP(n1207), .ZN(issueqPacket1_o[108]) );
  INVX0 U1218 ( .INP(renamedPacket1_i[108]), .ZN(n1207) );
  INVX0 U1219 ( .INP(n1209), .ZN(issueqPacket1_o[109]) );
  INVX0 U1220 ( .INP(renamedPacket1_i[109]), .ZN(n1209) );
  INVX0 U1221 ( .INP(n1211), .ZN(issueqPacket1_o[110]) );
  INVX0 U1222 ( .INP(renamedPacket1_i[110]), .ZN(n1211) );
  INVX0 U1223 ( .INP(n1213), .ZN(issueqPacket1_o[111]) );
  INVX0 U1224 ( .INP(renamedPacket1_i[111]), .ZN(n1213) );
  INVX0 U1225 ( .INP(n1215), .ZN(issueqPacket1_o[112]) );
  INVX0 U1226 ( .INP(renamedPacket1_i[112]), .ZN(n1215) );
  INVX0 U1227 ( .INP(n1217), .ZN(issueqPacket1_o[113]) );
  INVX0 U1228 ( .INP(renamedPacket1_i[113]), .ZN(n1217) );
  INVX0 U1229 ( .INP(n1243), .ZN(issueqPacket1_o[122]) );
  INVX0 U1230 ( .INP(renamedPacket1_i[122]), .ZN(n1243) );
  INVX0 U1231 ( .INP(n1266), .ZN(issueqPacket1_o[130]) );
  INVX0 U1232 ( .INP(renamedPacket1_i[130]), .ZN(n1266) );
  INVX0 U1233 ( .INP(n1268), .ZN(issueqPacket1_o[131]) );
  INVX0 U1234 ( .INP(renamedPacket1_i[131]), .ZN(n1268) );
  INVX0 U1235 ( .INP(n1278), .ZN(issueqPacket1_o[138]) );
  INVX0 U1236 ( .INP(issueqPacket1_o_138), .ZN(n1278) );
  INVX0 U1237 ( .INP(n1298), .ZN(issueqPacket0_o[0]) );
  INVX0 U1238 ( .INP(issueqPacket0_o_0), .ZN(n1298) );
  INVX0 U1239 ( .INP(n1300), .ZN(issueqPacket0_o[1]) );
  INVX0 U1240 ( .INP(issueqPacket0_o_1), .ZN(n1300) );
  INVX0 U1241 ( .INP(n1302), .ZN(issueqPacket0_o[2]) );
  INVX0 U1242 ( .INP(issueqPacket0_o_2), .ZN(n1302) );
  INVX0 U1243 ( .INP(n1304), .ZN(issueqPacket0_o[3]) );
  INVX0 U1244 ( .INP(issueqPacket0_o_3), .ZN(n1304) );
  INVX0 U1245 ( .INP(n1306), .ZN(issueqPacket0_o[4]) );
  INVX0 U1246 ( .INP(issueqPacket0_o_4), .ZN(n1306) );
  INVX0 U1247 ( .INP(n1308), .ZN(issueqPacket0_o[5]) );
  INVX0 U1248 ( .INP(issueqPacket0_o_5), .ZN(n1308) );
  INVX0 U1249 ( .INP(n1310), .ZN(issueqPacket0_o[6]) );
  INVX0 U1250 ( .INP(issueqPacket0_o_6), .ZN(n1310) );
  INVX0 U1251 ( .INP(n1312), .ZN(issueqPacket0_o[7]) );
  INVX0 U1252 ( .INP(issueqPacket0_o_7), .ZN(n1312) );
  INVX0 U1253 ( .INP(n1314), .ZN(issueqPacket0_o[8]) );
  INVX0 U1254 ( .INP(issueqPacket0_o_8), .ZN(n1314) );
  INVX0 U1255 ( .INP(n1316), .ZN(issueqPacket0_o[9]) );
  INVX0 U1256 ( .INP(issueqPacket0_o_9), .ZN(n1316) );
  INVX0 U1257 ( .INP(n1318), .ZN(issueqPacket0_o[10]) );
  INVX0 U1258 ( .INP(issueqPacket0_o_10), .ZN(n1318) );
  INVX0 U1259 ( .INP(n1320), .ZN(issueqPacket0_o[11]) );
  INVX0 U1260 ( .INP(issueqPacket0_o_11), .ZN(n1320) );
  INVX0 U1261 ( .INP(n1322), .ZN(issueqPacket0_o[12]) );
  INVX0 U1262 ( .INP(issueqPacket0_o_12), .ZN(n1322) );
  INVX0 U1263 ( .INP(n1324), .ZN(issueqPacket0_o[13]) );
  INVX0 U1264 ( .INP(issueqPacket0_o_13), .ZN(n1324) );
  INVX0 U1265 ( .INP(n1326), .ZN(issueqPacket0_o[14]) );
  INVX0 U1266 ( .INP(issueqPacket0_o_14), .ZN(n1326) );
  INVX0 U1267 ( .INP(n1328), .ZN(issueqPacket0_o[15]) );
  INVX0 U1268 ( .INP(issueqPacket0_o_15), .ZN(n1328) );
  INVX0 U1269 ( .INP(n1330), .ZN(issueqPacket0_o[16]) );
  INVX0 U1270 ( .INP(issueqPacket0_o_16), .ZN(n1330) );
  INVX0 U1271 ( .INP(n1332), .ZN(issueqPacket0_o[17]) );
  INVX0 U1272 ( .INP(issueqPacket0_o_17), .ZN(n1332) );
  INVX0 U1273 ( .INP(n1334), .ZN(issueqPacket0_o[18]) );
  INVX0 U1274 ( .INP(issueqPacket0_o_18), .ZN(n1334) );
  INVX0 U1275 ( .INP(n1336), .ZN(issueqPacket0_o[19]) );
  INVX0 U1276 ( .INP(issueqPacket0_o_19), .ZN(n1336) );
  INVX0 U1277 ( .INP(n1338), .ZN(issueqPacket0_o[20]) );
  INVX0 U1278 ( .INP(issueqPacket0_o_20), .ZN(n1338) );
  INVX0 U1279 ( .INP(n1340), .ZN(issueqPacket0_o[21]) );
  INVX0 U1280 ( .INP(issueqPacket0_o_21), .ZN(n1340) );
  INVX0 U1281 ( .INP(n1342), .ZN(issueqPacket0_o[22]) );
  INVX0 U1282 ( .INP(issueqPacket0_o_22), .ZN(n1342) );
  INVX0 U1283 ( .INP(n1344), .ZN(issueqPacket0_o[23]) );
  INVX0 U1284 ( .INP(issueqPacket0_o_23), .ZN(n1344) );
  INVX0 U1285 ( .INP(n1346), .ZN(issueqPacket0_o[24]) );
  INVX0 U1286 ( .INP(issueqPacket0_o_24), .ZN(n1346) );
  INVX0 U1287 ( .INP(n1348), .ZN(issueqPacket0_o[25]) );
  INVX0 U1288 ( .INP(issueqPacket0_o_25), .ZN(n1348) );
  INVX0 U1289 ( .INP(n1350), .ZN(issueqPacket0_o[26]) );
  INVX0 U1290 ( .INP(issueqPacket0_o_26), .ZN(n1350) );
  INVX0 U1291 ( .INP(n1352), .ZN(issueqPacket0_o[27]) );
  INVX0 U1292 ( .INP(issueqPacket0_o_27), .ZN(n1352) );
  INVX0 U1293 ( .INP(n1354), .ZN(issueqPacket0_o[28]) );
  INVX0 U1294 ( .INP(issueqPacket0_o_28), .ZN(n1354) );
  INVX0 U1295 ( .INP(n1356), .ZN(issueqPacket0_o[29]) );
  INVX0 U1296 ( .INP(issueqPacket0_o_29), .ZN(n1356) );
  INVX0 U1297 ( .INP(n1358), .ZN(issueqPacket0_o[30]) );
  INVX0 U1298 ( .INP(issueqPacket0_o_30), .ZN(n1358) );
  INVX0 U1299 ( .INP(n1360), .ZN(issueqPacket0_o[31]) );
  INVX0 U1300 ( .INP(issueqPacket0_o_31), .ZN(n1360) );
  INVX0 U1301 ( .INP(n1362), .ZN(issueqPacket0_o[32]) );
  INVX0 U1302 ( .INP(issueqPacket0_o_32), .ZN(n1362) );
  INVX0 U1303 ( .INP(n1364), .ZN(issueqPacket0_o[33]) );
  INVX0 U1304 ( .INP(issueqPacket0_o_33), .ZN(n1364) );
  INVX0 U1305 ( .INP(n1366), .ZN(issueqPacket0_o[34]) );
  INVX0 U1306 ( .INP(issueqPacket0_o_34), .ZN(n1366) );
  INVX0 U1307 ( .INP(n1368), .ZN(issueqPacket0_o[35]) );
  INVX0 U1308 ( .INP(issueqPacket0_o_35), .ZN(n1368) );
  INVX0 U1309 ( .INP(n1370), .ZN(issueqPacket0_o[36]) );
  INVX0 U1310 ( .INP(issueqPacket0_o_36), .ZN(n1370) );
  INVX0 U1311 ( .INP(n1372), .ZN(issueqPacket0_o[69]) );
  INVX0 U1312 ( .INP(renamedPacket0_i[69]), .ZN(n1372) );
  INVX0 U1313 ( .INP(n1374), .ZN(issueqPacket0_o[70]) );
  INVX0 U1314 ( .INP(renamedPacket0_i[70]), .ZN(n1374) );
  INVX0 U1315 ( .INP(n1376), .ZN(issueqPacket0_o[71]) );
  INVX0 U1316 ( .INP(renamedPacket0_i[71]), .ZN(n1376) );
  INVX0 U1317 ( .INP(n1378), .ZN(issueqPacket0_o[72]) );
  INVX0 U1318 ( .INP(renamedPacket0_i[72]), .ZN(n1378) );
  INVX0 U1319 ( .INP(n1380), .ZN(issueqPacket0_o[73]) );
  INVX0 U1320 ( .INP(renamedPacket0_i[73]), .ZN(n1380) );
  INVX0 U1321 ( .INP(n1382), .ZN(issueqPacket0_o[74]) );
  INVX0 U1322 ( .INP(renamedPacket0_i[74]), .ZN(n1382) );
  INVX0 U1323 ( .INP(n1384), .ZN(issueqPacket0_o[75]) );
  INVX0 U1324 ( .INP(renamedPacket0_i[75]), .ZN(n1384) );
  INVX0 U1325 ( .INP(n1386), .ZN(issueqPacket0_o[76]) );
  INVX0 U1326 ( .INP(renamedPacket0_i[76]), .ZN(n1386) );
  INVX0 U1327 ( .INP(n1388), .ZN(issueqPacket0_o[77]) );
  INVX0 U1328 ( .INP(renamedPacket0_i[77]), .ZN(n1388) );
  INVX0 U1329 ( .INP(n1390), .ZN(issueqPacket0_o[78]) );
  INVX0 U1330 ( .INP(renamedPacket0_i[78]), .ZN(n1390) );
  INVX0 U1331 ( .INP(n1392), .ZN(issueqPacket0_o[79]) );
  INVX0 U1332 ( .INP(renamedPacket0_i[79]), .ZN(n1392) );
  INVX0 U1333 ( .INP(n1394), .ZN(issueqPacket0_o[80]) );
  INVX0 U1334 ( .INP(renamedPacket0_i[80]), .ZN(n1394) );
  INVX0 U1335 ( .INP(n1396), .ZN(issueqPacket0_o[81]) );
  INVX0 U1336 ( .INP(renamedPacket0_i[81]), .ZN(n1396) );
  INVX0 U1337 ( .INP(n1398), .ZN(issueqPacket0_o[82]) );
  INVX0 U1338 ( .INP(renamedPacket0_i[82]), .ZN(n1398) );
  INVX0 U1339 ( .INP(n1400), .ZN(issueqPacket0_o[83]) );
  INVX0 U1340 ( .INP(renamedPacket0_i[83]), .ZN(n1400) );
  INVX0 U1341 ( .INP(n1402), .ZN(issueqPacket0_o[84]) );
  INVX0 U1342 ( .INP(renamedPacket0_i[84]), .ZN(n1402) );
  INVX0 U1343 ( .INP(n1404), .ZN(issueqPacket0_o[85]) );
  INVX0 U1344 ( .INP(renamedPacket0_i[85]), .ZN(n1404) );
  INVX0 U1345 ( .INP(n1406), .ZN(issueqPacket0_o[86]) );
  INVX0 U1346 ( .INP(renamedPacket0_i[86]), .ZN(n1406) );
  INVX0 U1347 ( .INP(n1408), .ZN(issueqPacket0_o[87]) );
  INVX0 U1348 ( .INP(renamedPacket0_i[87]), .ZN(n1408) );
  INVX0 U1349 ( .INP(n1410), .ZN(issueqPacket0_o[88]) );
  INVX0 U1350 ( .INP(renamedPacket0_i[88]), .ZN(n1410) );
  INVX0 U1351 ( .INP(n1412), .ZN(issueqPacket0_o[89]) );
  INVX0 U1352 ( .INP(renamedPacket0_i[89]), .ZN(n1412) );
  INVX0 U1353 ( .INP(n1414), .ZN(issueqPacket0_o[90]) );
  INVX0 U1354 ( .INP(renamedPacket0_i[90]), .ZN(n1414) );
  INVX0 U1355 ( .INP(n1416), .ZN(issueqPacket0_o[91]) );
  INVX0 U1356 ( .INP(renamedPacket0_i[91]), .ZN(n1416) );
  INVX0 U1357 ( .INP(n1418), .ZN(issueqPacket0_o[92]) );
  INVX0 U1358 ( .INP(renamedPacket0_i[92]), .ZN(n1418) );
  INVX0 U1359 ( .INP(n1420), .ZN(issueqPacket0_o[93]) );
  INVX0 U1360 ( .INP(renamedPacket0_i[93]), .ZN(n1420) );
  INVX0 U1361 ( .INP(n1422), .ZN(issueqPacket0_o[94]) );
  INVX0 U1362 ( .INP(renamedPacket0_i[94]), .ZN(n1422) );
  INVX0 U1363 ( .INP(n1424), .ZN(issueqPacket0_o[95]) );
  INVX0 U1364 ( .INP(renamedPacket0_i[95]), .ZN(n1424) );
  INVX0 U1365 ( .INP(n1426), .ZN(issueqPacket0_o[96]) );
  INVX0 U1366 ( .INP(renamedPacket0_i[96]), .ZN(n1426) );
  INVX0 U1367 ( .INP(n1428), .ZN(issueqPacket0_o[97]) );
  INVX0 U1368 ( .INP(renamedPacket0_i[97]), .ZN(n1428) );
  INVX0 U1369 ( .INP(n1430), .ZN(issueqPacket0_o[98]) );
  INVX0 U1370 ( .INP(renamedPacket0_i[98]), .ZN(n1430) );
  INVX0 U1371 ( .INP(n1432), .ZN(issueqPacket0_o[99]) );
  INVX0 U1372 ( .INP(renamedPacket0_i[99]), .ZN(n1432) );
  INVX0 U1373 ( .INP(n1434), .ZN(issueqPacket0_o[100]) );
  INVX0 U1374 ( .INP(renamedPacket0_i[100]), .ZN(n1434) );
  INVX0 U1375 ( .INP(n1436), .ZN(issueqPacket0_o[101]) );
  INVX0 U1376 ( .INP(renamedPacket0_i[101]), .ZN(n1436) );
  INVX0 U1377 ( .INP(n1438), .ZN(issueqPacket0_o[102]) );
  INVX0 U1378 ( .INP(renamedPacket0_i[102]), .ZN(n1438) );
  INVX0 U1379 ( .INP(n1440), .ZN(issueqPacket0_o[103]) );
  INVX0 U1380 ( .INP(renamedPacket0_i[103]), .ZN(n1440) );
  INVX0 U1381 ( .INP(n1442), .ZN(issueqPacket0_o[104]) );
  INVX0 U1382 ( .INP(renamedPacket0_i[104]), .ZN(n1442) );
  INVX0 U1383 ( .INP(n1444), .ZN(issueqPacket0_o[105]) );
  INVX0 U1384 ( .INP(renamedPacket0_i[105]), .ZN(n1444) );
  INVX0 U1385 ( .INP(n1446), .ZN(issueqPacket0_o[106]) );
  INVX0 U1386 ( .INP(renamedPacket0_i[106]), .ZN(n1446) );
  INVX0 U1387 ( .INP(n1448), .ZN(issueqPacket0_o[107]) );
  INVX0 U1388 ( .INP(renamedPacket0_i[107]), .ZN(n1448) );
  INVX0 U1389 ( .INP(n1450), .ZN(issueqPacket0_o[108]) );
  INVX0 U1390 ( .INP(renamedPacket0_i[108]), .ZN(n1450) );
  INVX0 U1391 ( .INP(n1452), .ZN(issueqPacket0_o[109]) );
  INVX0 U1392 ( .INP(renamedPacket0_i[109]), .ZN(n1452) );
  INVX0 U1393 ( .INP(n1454), .ZN(issueqPacket0_o[110]) );
  INVX0 U1394 ( .INP(renamedPacket0_i[110]), .ZN(n1454) );
  INVX0 U1395 ( .INP(n1456), .ZN(issueqPacket0_o[111]) );
  INVX0 U1396 ( .INP(renamedPacket0_i[111]), .ZN(n1456) );
  INVX0 U1397 ( .INP(n1458), .ZN(issueqPacket0_o[112]) );
  INVX0 U1398 ( .INP(renamedPacket0_i[112]), .ZN(n1458) );
  INVX0 U1399 ( .INP(n1460), .ZN(issueqPacket0_o[113]) );
  INVX0 U1400 ( .INP(renamedPacket0_i[113]), .ZN(n1460) );
  INVX0 U1401 ( .INP(n1462), .ZN(issueqPacket0_o[122]) );
  INVX0 U1402 ( .INP(issueqPacket0_o_122), .ZN(n1462) );
  INVX0 U1403 ( .INP(n1464), .ZN(issueqPacket0_o[130]) );
  INVX0 U1404 ( .INP(issueqPacket0_o_130), .ZN(n1464) );
  INVX0 U1405 ( .INP(n1466), .ZN(issueqPacket0_o[131]) );
  INVX0 U1406 ( .INP(issueqPacket0_o_131), .ZN(n1466) );
  INVX0 U1407 ( .INP(n1468), .ZN(issueqPacket0_o[138]) );
  INVX0 U1408 ( .INP(issueqPacket0_o_138), .ZN(n1468) );
  NAND2X1 U1409 ( .IN1(N9), .IN2(renamedPacket0_i[137]), .QN(n1480) );
  NAND2X1 U1410 ( .IN1(N4), .IN2(renamedPacket0_i[136]), .QN(n1482) );
  NOR2X0 U1411 ( .IN1(flagRecoverEX_i), .IN2(stallfrontEnd_o), .QN(n65) );
  INVX0 U1412 ( .INP(activeListCnt_i[2]), .ZN(N45) );
  INVX0 U1413 ( .INP(issueQueueCnt_i[2]), .ZN(N38) );
  INVX0 U1414 ( .INP(renamedPacket3_i[54]), .ZN(n414) );
  INVX0 U1415 ( .INP(renamedPacket3_i[55]), .ZN(n417) );
  INVX0 U1416 ( .INP(renamedPacket3_i[56]), .ZN(n420) );
  INVX0 U1417 ( .INP(renamedPacket3_i[57]), .ZN(n423) );
  INVX0 U1418 ( .INP(renamedPacket3_i[58]), .ZN(n426) );
  INVX0 U1419 ( .INP(renamedPacket3_i[59]), .ZN(n429) );
  INVX0 U1420 ( .INP(renamedPacket3_i[60]), .ZN(n432) );
  INVX0 U1421 ( .INP(renamedPacket3_i[61]), .ZN(n435) );
  INVX0 U1422 ( .INP(renamedPacket3_i[62]), .ZN(n438) );
  INVX0 U1423 ( .INP(renamedPacket3_i[63]), .ZN(n441) );
  INVX0 U1424 ( .INP(renamedPacket3_i[64]), .ZN(n444) );
  INVX0 U1425 ( .INP(renamedPacket3_i[65]), .ZN(n447) );
  INVX0 U1426 ( .INP(renamedPacket3_i[66]), .ZN(n450) );
  INVX0 U1427 ( .INP(renamedPacket3_i[67]), .ZN(n453) );
  INVX0 U1428 ( .INP(renamedPacket3_i[68]), .ZN(n456) );
  INVX0 U1429 ( .INP(renamedPacket3_i[69]), .ZN(n459) );
  INVX0 U1430 ( .INP(n459), .ZN(issueqPacket3_o[69]) );
  INVX0 U1431 ( .INP(n456), .ZN(issueqPacket3_o[68]) );
  INVX0 U1432 ( .INP(n456), .ZN(alPacket3_o[52]) );
  INVX0 U1433 ( .INP(n453), .ZN(issueqPacket3_o[67]) );
  INVX0 U1434 ( .INP(n453), .ZN(alPacket3_o[51]) );
  INVX0 U1435 ( .INP(n450), .ZN(issueqPacket3_o[66]) );
  INVX0 U1436 ( .INP(n450), .ZN(alPacket3_o[50]) );
  INVX0 U1437 ( .INP(n447), .ZN(issueqPacket3_o[65]) );
  INVX0 U1438 ( .INP(n447), .ZN(alPacket3_o[49]) );
  INVX0 U1439 ( .INP(n444), .ZN(issueqPacket3_o[64]) );
  INVX0 U1440 ( .INP(n444), .ZN(alPacket3_o[48]) );
  INVX0 U1441 ( .INP(n441), .ZN(issueqPacket3_o[63]) );
  INVX0 U1442 ( .INP(n441), .ZN(alPacket3_o[47]) );
  INVX0 U1443 ( .INP(n438), .ZN(issueqPacket3_o[62]) );
  INVX0 U1444 ( .INP(n438), .ZN(alPacket3_o[46]) );
  INVX0 U1445 ( .INP(n435), .ZN(issueqPacket3_o[61]) );
  INVX0 U1446 ( .INP(n435), .ZN(alPacket3_o[45]) );
  INVX0 U1447 ( .INP(n432), .ZN(issueqPacket3_o[60]) );
  INVX0 U1448 ( .INP(n432), .ZN(alPacket3_o[44]) );
  INVX0 U1449 ( .INP(n429), .ZN(issueqPacket3_o[59]) );
  INVX0 U1450 ( .INP(n429), .ZN(alPacket3_o[43]) );
  INVX0 U1451 ( .INP(n426), .ZN(issueqPacket3_o[58]) );
  INVX0 U1452 ( .INP(n426), .ZN(alPacket3_o[42]) );
  INVX0 U1453 ( .INP(n423), .ZN(issueqPacket3_o[57]) );
  INVX0 U1454 ( .INP(n423), .ZN(alPacket3_o[41]) );
  INVX0 U1455 ( .INP(n420), .ZN(issueqPacket3_o[56]) );
  INVX0 U1456 ( .INP(n420), .ZN(alPacket3_o[40]) );
  INVX0 U1457 ( .INP(n417), .ZN(issueqPacket3_o[55]) );
  INVX0 U1458 ( .INP(n417), .ZN(alPacket3_o[39]) );
  INVX0 U1459 ( .INP(n414), .ZN(issueqPacket3_o[54]) );
  INVX0 U1460 ( .INP(n414), .ZN(alPacket3_o[38]) );
  AND2X1 U1461 ( .IN1(issueQueueCnt_i[5]), .IN2(\add_290/carry[5] ), .Q(N42)
         );
  XOR2X1 U1462 ( .IN1(\add_290/carry[5] ), .IN2(issueQueueCnt_i[5]), .Q(N41)
         );
  AND2X1 U1463 ( .IN1(issueQueueCnt_i[4]), .IN2(\add_290/carry[4] ), .Q(
        \add_290/carry[5] ) );
  XOR2X1 U1464 ( .IN1(\add_290/carry[4] ), .IN2(issueQueueCnt_i[4]), .Q(N40)
         );
  AND2X1 U1465 ( .IN1(issueQueueCnt_i[3]), .IN2(issueQueueCnt_i[2]), .Q(
        \add_290/carry[4] ) );
  XOR2X1 U1466 ( .IN1(issueQueueCnt_i[2]), .IN2(issueQueueCnt_i[3]), .Q(N39)
         );
  AND2X1 U1467 ( .IN1(activeListCnt_i[7]), .IN2(\add_291/carry[7] ), .Q(N51)
         );
  XOR2X1 U1468 ( .IN1(\add_291/carry[7] ), .IN2(activeListCnt_i[7]), .Q(N50)
         );
  AND2X1 U1469 ( .IN1(activeListCnt_i[6]), .IN2(\add_291/carry[6] ), .Q(
        \add_291/carry[7] ) );
  XOR2X1 U1470 ( .IN1(\add_291/carry[6] ), .IN2(activeListCnt_i[6]), .Q(N49)
         );
  AND2X1 U1471 ( .IN1(activeListCnt_i[5]), .IN2(\add_291/carry[5] ), .Q(
        \add_291/carry[6] ) );
  XOR2X1 U1472 ( .IN1(\add_291/carry[5] ), .IN2(activeListCnt_i[5]), .Q(N48)
         );
  AND2X1 U1473 ( .IN1(activeListCnt_i[4]), .IN2(\add_291/carry[4] ), .Q(
        \add_291/carry[5] ) );
  XOR2X1 U1474 ( .IN1(\add_291/carry[4] ), .IN2(activeListCnt_i[4]), .Q(N47)
         );
  AND2X1 U1475 ( .IN1(activeListCnt_i[3]), .IN2(activeListCnt_i[2]), .Q(
        \add_291/carry[4] ) );
  XOR2X1 U1476 ( .IN1(activeListCnt_i[2]), .IN2(activeListCnt_i[3]), .Q(N46)
         );
  AND2X1 U1477 ( .IN1(loadQueueCnt_i[5]), .IN2(\add_288/carry[5] ), .Q(N28) );
  XOR2X1 U1478 ( .IN1(\add_288/carry[5] ), .IN2(loadQueueCnt_i[5]), .Q(N27) );
  AND2X1 U1479 ( .IN1(loadQueueCnt_i[4]), .IN2(\add_288/carry[4] ), .Q(
        \add_288/carry[5] ) );
  XOR2X1 U1480 ( .IN1(\add_288/carry[4] ), .IN2(loadQueueCnt_i[4]), .Q(N26) );
  AND2X1 U1481 ( .IN1(loadQueueCnt_i[3]), .IN2(\add_288/carry[3] ), .Q(
        \add_288/carry[4] ) );
  XOR2X1 U1482 ( .IN1(\add_288/carry[3] ), .IN2(loadQueueCnt_i[3]), .Q(N25) );
  AND2X1 U1483 ( .IN1(loadQueueCnt_i[0]), .IN2(\loadCnt[0] ), .Q(
        \add_288/carry[1] ) );
  XOR2X1 U1484 ( .IN1(\loadCnt[0] ), .IN2(loadQueueCnt_i[0]), .Q(N22) );
  AND2X1 U1485 ( .IN1(storeQueueCnt_i[5]), .IN2(\add_289/carry[5] ), .Q(N35)
         );
  XOR2X1 U1486 ( .IN1(\add_289/carry[5] ), .IN2(storeQueueCnt_i[5]), .Q(N34)
         );
  AND2X1 U1487 ( .IN1(storeQueueCnt_i[4]), .IN2(\add_289/carry[4] ), .Q(
        \add_289/carry[5] ) );
  XOR2X1 U1488 ( .IN1(\add_289/carry[4] ), .IN2(storeQueueCnt_i[4]), .Q(N33)
         );
  AND2X1 U1489 ( .IN1(storeQueueCnt_i[3]), .IN2(\add_289/carry[3] ), .Q(
        \add_289/carry[4] ) );
  XOR2X1 U1490 ( .IN1(\add_289/carry[3] ), .IN2(storeQueueCnt_i[3]), .Q(N32)
         );
  AND2X1 U1491 ( .IN1(storeQueueCnt_i[0]), .IN2(\storeCnt[0] ), .Q(
        \add_289/carry[1] ) );
  XOR2X1 U1492 ( .IN1(\storeCnt[0] ), .IN2(storeQueueCnt_i[0]), .Q(N29) );
  OR3X1 U1493 ( .IN1(N28), .IN2(N26), .IN3(N25), .Q(n1470) );
  OR4X1 U1494 ( .IN1(N24), .IN2(N23), .IN3(N22), .IN4(n1470), .Q(n1471) );
  OA21X1 U1495 ( .IN1(N28), .IN2(N27), .IN3(n1471), .Q(stall0) );
  OR3X1 U1496 ( .IN1(N35), .IN2(N33), .IN3(N32), .Q(n1472) );
  OR4X1 U1497 ( .IN1(N31), .IN2(N30), .IN3(N29), .IN4(n1472), .Q(n1473) );
  OA21X1 U1498 ( .IN1(N35), .IN2(N34), .IN3(n1473), .Q(stall1) );
  OR3X1 U1499 ( .IN1(N42), .IN2(N40), .IN3(N39), .Q(n1474) );
  OR4X1 U1500 ( .IN1(N38), .IN2(N37), .IN3(N36), .IN4(n1474), .Q(n1475) );
  OA21X1 U1501 ( .IN1(N42), .IN2(N41), .IN3(n1475), .Q(stall2) );
  OR4X1 U1502 ( .IN1(N47), .IN2(N46), .IN3(N49), .IN4(N48), .Q(n1476) );
  OR4X1 U1503 ( .IN1(N45), .IN2(N44), .IN3(N43), .IN4(n1476), .Q(n1477) );
  AO21X1 U1504 ( .IN1(N50), .IN2(n1477), .IN3(N51), .Q(stall3) );
  AND3X1 U1505 ( .IN1(N10), .IN2(renamedPacket0_i[137]), .IN3(N9), .Q(
        \storeCnt[2] ) );
  XNOR2X1 U1506 ( .IN1(N10), .IN2(n1480), .Q(\storeCnt[1] ) );
  XOR2X1 U1507 ( .IN1(N9), .IN2(renamedPacket0_i[137]), .Q(\storeCnt[0] ) );
  AO22X1 U1508 ( .IN1(issueqPacket2_o_137), .IN2(issueqPacket1_o_137), .IN3(
        renamedPacket3_i[137]), .IN4(n1481), .Q(N10) );
  XOR2X1 U1509 ( .IN1(renamedPacket3_i[137]), .IN2(n1481), .Q(N9) );
  XOR2X1 U1510 ( .IN1(issueqPacket2_o_137), .IN2(issueqPacket1_o_137), .Q(
        n1481) );
  AND3X1 U1511 ( .IN1(N5), .IN2(renamedPacket0_i[136]), .IN3(N4), .Q(
        \loadCnt[2] ) );
  XNOR2X1 U1512 ( .IN1(N5), .IN2(n1482), .Q(\loadCnt[1] ) );
  XOR2X1 U1513 ( .IN1(N4), .IN2(renamedPacket0_i[136]), .Q(\loadCnt[0] ) );
  AO22X1 U1514 ( .IN1(issueqPacket2_o_136), .IN2(issueqPacket1_o_136), .IN3(
        renamedPacket3_i[136]), .IN4(n1483), .Q(N5) );
  XOR2X1 U1515 ( .IN1(renamedPacket3_i[136]), .IN2(n1483), .Q(N4) );
  XOR2X1 U1516 ( .IN1(issueqPacket2_o_136), .IN2(issueqPacket1_o_136), .Q(
        n1483) );
endmodule

