
module WriteBack ( exePacketValid0_i, exePacket0_i, writebkValid0_o, ctrlFU0_o, 
        bypassValid0_o, bypassPacket0_o, computedAddr0_o, exePacketValid1_i, 
        exePacket1_i, writebkValid1_o, ctrlFU1_o, bypassValid1_o, 
        bypassPacket1_o, computedAddr1_o, exePacketValid2_i, exePacket2_i, 
        writebkValid2_o, ctrlFU2_o, bypassValid2_o, bypassPacket2_o, 
        computedAddr2_o, exePacketValid3_i, exePacket3_i, writebkValid3_o, 
        ctrlFU3_o, bypassValid3_o, bypassPacket3_o, computedAddr3_o, 
        lsuPacketValid0_i, lsuPacket0_i, ldViolationPacket_i, 
        agenIqFreedValid0_o, agenIqEntry0_o, ctrlVerified_o, ctrlMispredict_o, 
        ctrlConditional_o, ctrlSMTid_o, ctrlTargetAddr_o, ctrlBrDirection_o, 
        ctrlCtiQueueIndex_o, ldViolationPacket_o, clk, reset );
  input [106:0] exePacket0_i;
  output [14:0] ctrlFU0_o;
  output [41:0] bypassPacket0_o;
  output [31:0] computedAddr0_o;
  input [106:0] exePacket1_i;
  output [14:0] ctrlFU1_o;
  output [41:0] bypassPacket1_o;
  output [31:0] computedAddr1_o;
  input [106:0] exePacket2_i;
  output [14:0] ctrlFU2_o;
  output [41:0] bypassPacket2_o;
  output [31:0] computedAddr2_o;
  input [108:0] exePacket3_i;
  output [14:0] ctrlFU3_o;
  output [41:0] bypassPacket3_o;
  output [31:0] computedAddr3_o;
  input [62:0] lsuPacket0_i;
  input [7:0] ldViolationPacket_i;
  output [4:0] agenIqEntry0_o;
  output [1:0] ctrlSMTid_o;
  output [31:0] ctrlTargetAddr_o;
  output [3:0] ctrlCtiQueueIndex_o;
  output [7:0] ldViolationPacket_o;
  input exePacketValid0_i, exePacketValid1_i, exePacketValid2_i,
         exePacketValid3_i, lsuPacketValid0_i, clk, reset;
  output writebkValid0_o, bypassValid0_o, writebkValid1_o, bypassValid1_o,
         writebkValid2_o, bypassValid2_o, writebkValid3_o, bypassValid3_o,
         agenIqFreedValid0_o, ctrlVerified_o, ctrlMispredict_o,
         ctrlConditional_o, ctrlBrDirection_o;
  wire   exePacket0_i_38, exePacket0_i_37, exePacket1_i_38, exePacket1_i_37,
         exePacket2_i_38, exePacket2_i_37, exePacket2_i_36, exePacket2_i_35,
         exePacket2_i_34, exePacket2_i_33, exePacket2_i_32, exePacket2_i_31,
         exePacket2_i_30, exePacket2_i_29, exePacket2_i_28, exePacket2_i_27,
         exePacket2_i_26, exePacket2_i_25, exePacket2_i_24, exePacket2_i_23,
         exePacket2_i_22, exePacket2_i_21, exePacket2_i_20, exePacket2_i_19,
         exePacket2_i_18, exePacket2_i_17, exePacket2_i_16, exePacket2_i_15,
         exePacket2_i_14, exePacket2_i_13, exePacket2_i_12, exePacket2_i_11,
         exePacket2_i_10, exePacket2_i_9, exePacket2_i_8, exePacket2_i_7,
         exePacket2_i_6, exePacket2_i_5, exePacket2_i_4, exePacket2_i_3,
         exePacket2_i_2, exePacket2_i_1, exePacket2_i_0, exePacketValid0,
         exePacketValid1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n561, n563, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593;
  assign exePacket0_i_38 = exePacket0_i[38];
  assign exePacket0_i_37 = exePacket0_i[37];
  assign exePacket1_i_38 = exePacket1_i[38];
  assign exePacket1_i_37 = exePacket1_i[37];
  assign exePacket2_i_38 = exePacket2_i[38];
  assign exePacket2_i_37 = exePacket2_i[37];
  assign exePacket2_i_36 = exePacket2_i[36];
  assign exePacket2_i_35 = exePacket2_i[35];
  assign exePacket2_i_34 = exePacket2_i[34];
  assign exePacket2_i_33 = exePacket2_i[33];
  assign exePacket2_i_32 = exePacket2_i[32];
  assign exePacket2_i_31 = exePacket2_i[31];
  assign exePacket2_i_30 = exePacket2_i[30];
  assign exePacket2_i_29 = exePacket2_i[29];
  assign exePacket2_i_28 = exePacket2_i[28];
  assign exePacket2_i_27 = exePacket2_i[27];
  assign exePacket2_i_26 = exePacket2_i[26];
  assign exePacket2_i_25 = exePacket2_i[25];
  assign exePacket2_i_24 = exePacket2_i[24];
  assign exePacket2_i_23 = exePacket2_i[23];
  assign exePacket2_i_22 = exePacket2_i[22];
  assign exePacket2_i_21 = exePacket2_i[21];
  assign exePacket2_i_20 = exePacket2_i[20];
  assign exePacket2_i_19 = exePacket2_i[19];
  assign exePacket2_i_18 = exePacket2_i[18];
  assign exePacket2_i_17 = exePacket2_i[17];
  assign exePacket2_i_16 = exePacket2_i[16];
  assign exePacket2_i_15 = exePacket2_i[15];
  assign exePacket2_i_14 = exePacket2_i[14];
  assign exePacket2_i_13 = exePacket2_i[13];
  assign exePacket2_i_12 = exePacket2_i[12];
  assign exePacket2_i_11 = exePacket2_i[11];
  assign exePacket2_i_10 = exePacket2_i[10];
  assign exePacket2_i_9 = exePacket2_i[9];
  assign exePacket2_i_8 = exePacket2_i[8];
  assign exePacket2_i_7 = exePacket2_i[7];
  assign exePacket2_i_6 = exePacket2_i[6];
  assign exePacket2_i_5 = exePacket2_i[5];
  assign exePacket2_i_4 = exePacket2_i[4];
  assign exePacket2_i_3 = exePacket2_i[3];
  assign exePacket2_i_2 = exePacket2_i[2];
  assign exePacket2_i_1 = exePacket2_i[1];
  assign exePacket2_i_0 = exePacket2_i[0];
  assign writebkValid0_o = exePacketValid0;
  assign writebkValid1_o = exePacketValid1;

  DFFSSRX1 exePacketValid1_reg ( .D(n6), .RSTB(exePacketValid1_i), .SETB(1'b1), 
        .CLK(clk), .Q(exePacketValid1) );
  DFFSSRX1 lsuPacketValid0_reg ( .D(lsuPacketValid0_i), .RSTB(n6), .SETB(1'b1), 
        .CLK(clk), .Q(agenIqFreedValid0_o), .QN(n563) );
  DFFX1 \lsuPacket0_reg[58]  ( .D(n287), .CLK(clk), .Q(ctrlFU3_o[7]) );
  DFFX1 \lsuPacket0_reg[57]  ( .D(n286), .CLK(clk), .Q(ctrlFU3_o[6]) );
  DFFX1 \lsuPacket0_reg[56]  ( .D(n285), .CLK(clk), .Q(ctrlFU3_o[5]) );
  DFFX1 \lsuPacket0_reg[55]  ( .D(n284), .CLK(clk), .Q(ctrlFU3_o[4]) );
  DFFX1 \lsuPacket0_reg[54]  ( .D(n283), .CLK(clk), .Q(ctrlFU3_o[3]) );
  DFFX1 \lsuPacket0_reg[53]  ( .D(n282), .CLK(clk), .Q(ctrlFU3_o[2]) );
  DFFX1 \lsuPacket0_reg[52]  ( .D(n281), .CLK(clk), .Q(ctrlFU3_o[1]) );
  DFFX1 \lsuPacket0_reg[51]  ( .D(n280), .CLK(clk), .Q(ctrlFU3_o[0]) );
  DFFX1 \lsuPacket0_reg[50]  ( .D(n279), .CLK(clk), .Q(bypassPacket3_o[34]) );
  DFFX1 \lsuPacket0_reg[49]  ( .D(n278), .CLK(clk), .Q(bypassPacket3_o[33]) );
  DFFX1 \lsuPacket0_reg[48]  ( .D(n277), .CLK(clk), .Q(bypassPacket3_o[32]) );
  DFFX1 \lsuPacket0_reg[47]  ( .D(n276), .CLK(clk), .Q(bypassPacket3_o[31]) );
  DFFX1 \lsuPacket0_reg[46]  ( .D(n275), .CLK(clk), .Q(bypassPacket3_o[30]) );
  DFFX1 \lsuPacket0_reg[45]  ( .D(n274), .CLK(clk), .Q(bypassPacket3_o[29]) );
  DFFX1 \lsuPacket0_reg[44]  ( .D(n273), .CLK(clk), .Q(bypassPacket3_o[28]) );
  DFFX1 \lsuPacket0_reg[43]  ( .D(n272), .CLK(clk), .Q(bypassPacket3_o[27]) );
  DFFX1 \lsuPacket0_reg[42]  ( .D(n271), .CLK(clk), .Q(bypassPacket3_o[26]) );
  DFFX1 \lsuPacket0_reg[41]  ( .D(n270), .CLK(clk), .Q(bypassPacket3_o[25]) );
  DFFX1 \lsuPacket0_reg[40]  ( .D(n269), .CLK(clk), .Q(bypassPacket3_o[24]) );
  DFFX1 \lsuPacket0_reg[39]  ( .D(n268), .CLK(clk), .Q(bypassPacket3_o[23]) );
  DFFX1 \lsuPacket0_reg[38]  ( .D(n267), .CLK(clk), .Q(bypassPacket3_o[22]) );
  DFFX1 \lsuPacket0_reg[37]  ( .D(n266), .CLK(clk), .Q(bypassPacket3_o[21]) );
  DFFX1 \lsuPacket0_reg[36]  ( .D(n265), .CLK(clk), .Q(bypassPacket3_o[20]) );
  DFFX1 \lsuPacket0_reg[35]  ( .D(n264), .CLK(clk), .Q(bypassPacket3_o[19]) );
  DFFX1 \lsuPacket0_reg[34]  ( .D(n263), .CLK(clk), .Q(bypassPacket3_o[18]) );
  DFFX1 \lsuPacket0_reg[33]  ( .D(n262), .CLK(clk), .Q(bypassPacket3_o[17]) );
  DFFX1 \lsuPacket0_reg[32]  ( .D(n261), .CLK(clk), .Q(bypassPacket3_o[16]) );
  DFFX1 \lsuPacket0_reg[31]  ( .D(n260), .CLK(clk), .Q(bypassPacket3_o[15]) );
  DFFX1 \lsuPacket0_reg[30]  ( .D(n259), .CLK(clk), .Q(bypassPacket3_o[14]) );
  DFFX1 \lsuPacket0_reg[29]  ( .D(n258), .CLK(clk), .Q(bypassPacket3_o[13]) );
  DFFX1 \lsuPacket0_reg[28]  ( .D(n257), .CLK(clk), .Q(bypassPacket3_o[12]) );
  DFFX1 \lsuPacket0_reg[27]  ( .D(n256), .CLK(clk), .Q(bypassPacket3_o[11]) );
  DFFX1 \lsuPacket0_reg[26]  ( .D(n255), .CLK(clk), .Q(bypassPacket3_o[10]) );
  DFFX1 \lsuPacket0_reg[25]  ( .D(n254), .CLK(clk), .Q(bypassPacket3_o[9]) );
  DFFX1 \lsuPacket0_reg[24]  ( .D(n253), .CLK(clk), .Q(bypassPacket3_o[8]) );
  DFFX1 \lsuPacket0_reg[23]  ( .D(n252), .CLK(clk), .Q(bypassPacket3_o[7]) );
  DFFX1 \lsuPacket0_reg[22]  ( .D(n251), .CLK(clk), .Q(bypassPacket3_o[6]) );
  DFFX1 \lsuPacket0_reg[21]  ( .D(n250), .CLK(clk), .Q(bypassPacket3_o[5]) );
  DFFX1 \lsuPacket0_reg[20]  ( .D(n249), .CLK(clk), .Q(bypassPacket3_o[4]) );
  DFFX1 \lsuPacket0_reg[19]  ( .D(n248), .CLK(clk), .Q(bypassPacket3_o[3]) );
  DFFX1 \lsuPacket0_reg[18]  ( .D(n247), .CLK(clk), .Q(bypassPacket3_o[41]) );
  DFFX1 \lsuPacket0_reg[17]  ( .D(n246), .CLK(clk), .Q(bypassPacket3_o[40]) );
  DFFX1 \lsuPacket0_reg[16]  ( .D(n245), .CLK(clk), .Q(bypassPacket3_o[39]) );
  DFFX1 \lsuPacket0_reg[15]  ( .D(n244), .CLK(clk), .Q(bypassPacket3_o[38]) );
  DFFX1 \lsuPacket0_reg[14]  ( .D(n243), .CLK(clk), .Q(bypassPacket3_o[37]) );
  DFFX1 \lsuPacket0_reg[13]  ( .D(n242), .CLK(clk), .Q(bypassPacket3_o[36]) );
  DFFX1 \lsuPacket0_reg[12]  ( .D(n241), .CLK(clk), .Q(bypassPacket3_o[35]) );
  DFFX1 \lsuPacket0_reg[11]  ( .D(n240), .CLK(clk), .Q(ctrlFU3_o[14]) );
  DFFX1 \lsuPacket0_reg[10]  ( .D(n239), .CLK(clk), .Q(ctrlFU3_o[13]) );
  DFFX1 \lsuPacket0_reg[9]  ( .D(n238), .CLK(clk), .Q(ctrlFU3_o[12]) );
  DFFX1 \lsuPacket0_reg[8]  ( .D(n237), .CLK(clk), .Q(ctrlFU3_o[11]) );
  DFFX1 \lsuPacket0_reg[7]  ( .D(n236), .CLK(clk), .Q(ctrlFU3_o[10]) );
  DFFX1 \lsuPacket0_reg[6]  ( .D(n235), .CLK(clk), .Q(ctrlFU3_o[9]) );
  DFFX1 \lsuPacket0_reg[5]  ( .D(n234), .CLK(clk), .Q(ctrlFU3_o[8]) );
  DFFX1 \lsuPacket0_reg[4]  ( .D(n233), .CLK(clk), .Q(agenIqEntry0_o[4]) );
  DFFX1 \lsuPacket0_reg[3]  ( .D(n232), .CLK(clk), .Q(agenIqEntry0_o[3]) );
  DFFX1 \lsuPacket0_reg[2]  ( .D(n231), .CLK(clk), .Q(agenIqEntry0_o[2]) );
  DFFX1 \lsuPacket0_reg[1]  ( .D(n230), .CLK(clk), .Q(agenIqEntry0_o[1]) );
  DFFX1 \lsuPacket0_reg[0]  ( .D(n229), .CLK(clk), .Q(agenIqEntry0_o[0]) );
  DFFSSRX1 exePacketValid2_reg ( .D(n6), .RSTB(exePacketValid2_i), .SETB(1'b1), 
        .CLK(clk), .Q(ctrlVerified_o), .QN(n561) );
  DFFX1 \exePacket2_reg[102]  ( .D(n228), .CLK(clk), .Q(ctrlFU2_o[7]) );
  DFFX1 \exePacket2_reg[101]  ( .D(n227), .CLK(clk), .Q(ctrlFU2_o[6]) );
  DFFX1 \exePacket2_reg[100]  ( .D(n226), .CLK(clk), .Q(ctrlFU2_o[5]), .QN(
        n528) );
  DFFX1 \exePacket2_reg[99]  ( .D(n225), .CLK(clk), .Q(ctrlFU2_o[4]) );
  DFFX1 \exePacket2_reg[98]  ( .D(n224), .CLK(clk), .Q(ctrlFU2_o[3]) );
  DFFX1 \exePacket2_reg[97]  ( .D(n223), .CLK(clk), .Q(ctrlFU2_o[2]) );
  DFFX1 \exePacket2_reg[96]  ( .D(n222), .CLK(clk), .Q(ctrlFU2_o[1]) );
  DFFX1 \exePacket2_reg[95]  ( .D(n221), .CLK(clk), .Q(ctrlFU2_o[0]) );
  DFFX1 \exePacket2_reg[94]  ( .D(n220), .CLK(clk), .Q(bypassPacket2_o[41]) );
  DFFX1 \exePacket2_reg[93]  ( .D(n219), .CLK(clk), .Q(bypassPacket2_o[40]) );
  DFFX1 \exePacket2_reg[92]  ( .D(n218), .CLK(clk), .Q(bypassPacket2_o[39]) );
  DFFX1 \exePacket2_reg[91]  ( .D(n217), .CLK(clk), .Q(bypassPacket2_o[38]) );
  DFFX1 \exePacket2_reg[90]  ( .D(n216), .CLK(clk), .Q(bypassPacket2_o[37]) );
  DFFX1 \exePacket2_reg[89]  ( .D(n215), .CLK(clk), .Q(bypassPacket2_o[36]) );
  DFFX1 \exePacket2_reg[88]  ( .D(n214), .CLK(clk), .Q(bypassPacket2_o[35]) );
  DFFX1 \exePacket2_reg[87]  ( .D(n213), .CLK(clk), .Q(ctrlFU2_o[14]) );
  DFFX1 \exePacket2_reg[86]  ( .D(n212), .CLK(clk), .Q(ctrlFU2_o[13]) );
  DFFX1 \exePacket2_reg[85]  ( .D(n211), .CLK(clk), .Q(ctrlFU2_o[12]) );
  DFFX1 \exePacket2_reg[84]  ( .D(n210), .CLK(clk), .Q(ctrlFU2_o[11]) );
  DFFX1 \exePacket2_reg[83]  ( .D(n209), .CLK(clk), .Q(ctrlFU2_o[10]) );
  DFFX1 \exePacket2_reg[82]  ( .D(n208), .CLK(clk), .Q(ctrlFU2_o[9]) );
  DFFX1 \exePacket2_reg[81]  ( .D(n207), .CLK(clk), .Q(ctrlFU2_o[8]) );
  DFFX1 \exePacket2_reg[80]  ( .D(n206), .CLK(clk), .Q(bypassPacket2_o[34]) );
  DFFX1 \exePacket2_reg[79]  ( .D(n205), .CLK(clk), .Q(bypassPacket2_o[33]) );
  DFFX1 \exePacket2_reg[78]  ( .D(n204), .CLK(clk), .Q(bypassPacket2_o[32]) );
  DFFX1 \exePacket2_reg[77]  ( .D(n203), .CLK(clk), .Q(bypassPacket2_o[31]) );
  DFFX1 \exePacket2_reg[76]  ( .D(n202), .CLK(clk), .Q(bypassPacket2_o[30]) );
  DFFX1 \exePacket2_reg[75]  ( .D(n201), .CLK(clk), .Q(bypassPacket2_o[29]) );
  DFFX1 \exePacket2_reg[74]  ( .D(n200), .CLK(clk), .Q(bypassPacket2_o[28]) );
  DFFX1 \exePacket2_reg[73]  ( .D(n199), .CLK(clk), .Q(bypassPacket2_o[27]) );
  DFFX1 \exePacket2_reg[72]  ( .D(n198), .CLK(clk), .Q(bypassPacket2_o[26]) );
  DFFX1 \exePacket2_reg[71]  ( .D(n197), .CLK(clk), .Q(bypassPacket2_o[25]) );
  DFFX1 \exePacket2_reg[70]  ( .D(n196), .CLK(clk), .Q(bypassPacket2_o[24]) );
  DFFX1 \exePacket2_reg[69]  ( .D(n195), .CLK(clk), .Q(bypassPacket2_o[23]) );
  DFFX1 \exePacket2_reg[68]  ( .D(n194), .CLK(clk), .Q(bypassPacket2_o[22]) );
  DFFX1 \exePacket2_reg[67]  ( .D(n193), .CLK(clk), .Q(bypassPacket2_o[21]) );
  DFFX1 \exePacket2_reg[66]  ( .D(n192), .CLK(clk), .Q(bypassPacket2_o[20]) );
  DFFX1 \exePacket2_reg[65]  ( .D(n191), .CLK(clk), .Q(bypassPacket2_o[19]) );
  DFFX1 \exePacket2_reg[64]  ( .D(n190), .CLK(clk), .Q(bypassPacket2_o[18]) );
  DFFX1 \exePacket2_reg[63]  ( .D(n189), .CLK(clk), .Q(bypassPacket2_o[17]) );
  DFFX1 \exePacket2_reg[62]  ( .D(n188), .CLK(clk), .Q(bypassPacket2_o[16]) );
  DFFX1 \exePacket2_reg[61]  ( .D(n187), .CLK(clk), .Q(bypassPacket2_o[15]) );
  DFFX1 \exePacket2_reg[60]  ( .D(n186), .CLK(clk), .Q(bypassPacket2_o[14]) );
  DFFX1 \exePacket2_reg[59]  ( .D(n185), .CLK(clk), .Q(bypassPacket2_o[13]) );
  DFFX1 \exePacket2_reg[58]  ( .D(n184), .CLK(clk), .Q(bypassPacket2_o[12]) );
  DFFX1 \exePacket2_reg[57]  ( .D(n183), .CLK(clk), .Q(bypassPacket2_o[11]) );
  DFFX1 \exePacket2_reg[56]  ( .D(n182), .CLK(clk), .Q(bypassPacket2_o[10]) );
  DFFX1 \exePacket2_reg[55]  ( .D(n181), .CLK(clk), .Q(bypassPacket2_o[9]) );
  DFFX1 \exePacket2_reg[54]  ( .D(n180), .CLK(clk), .Q(bypassPacket2_o[8]) );
  DFFX1 \exePacket2_reg[53]  ( .D(n179), .CLK(clk), .Q(bypassPacket2_o[7]) );
  DFFX1 \exePacket2_reg[52]  ( .D(n178), .CLK(clk), .Q(bypassPacket2_o[6]) );
  DFFX1 \exePacket2_reg[51]  ( .D(n177), .CLK(clk), .Q(bypassPacket2_o[5]) );
  DFFX1 \exePacket2_reg[50]  ( .D(n176), .CLK(clk), .Q(bypassPacket2_o[4]) );
  DFFX1 \exePacket2_reg[49]  ( .D(n175), .CLK(clk), .Q(bypassPacket2_o[3]) );
  DFFX1 \exePacket2_reg[38]  ( .D(n174), .CLK(clk), .Q(bypassPacket2_o[2]), 
        .QN(n527) );
  DFFX1 \exePacket2_reg[37]  ( .D(n173), .CLK(clk), .Q(bypassPacket2_o[1]), 
        .QN(n526) );
  DFFX1 \exePacket2_reg[36]  ( .D(n172), .CLK(clk), .Q(ctrlCtiQueueIndex_o[3])
         );
  DFFX1 \exePacket2_reg[35]  ( .D(n171), .CLK(clk), .Q(ctrlCtiQueueIndex_o[2])
         );
  DFFX1 \exePacket2_reg[34]  ( .D(n170), .CLK(clk), .Q(ctrlCtiQueueIndex_o[1])
         );
  DFFX1 \exePacket2_reg[33]  ( .D(n169), .CLK(clk), .Q(ctrlCtiQueueIndex_o[0])
         );
  DFFX1 \exePacket2_reg[32]  ( .D(n168), .CLK(clk), .Q(computedAddr2_o[31]), 
        .QN(n525) );
  DFFX1 \exePacket2_reg[31]  ( .D(n167), .CLK(clk), .Q(computedAddr2_o[30]), 
        .QN(n524) );
  DFFX1 \exePacket2_reg[30]  ( .D(n166), .CLK(clk), .Q(computedAddr2_o[29]), 
        .QN(n523) );
  DFFX1 \exePacket2_reg[29]  ( .D(n165), .CLK(clk), .Q(computedAddr2_o[28]), 
        .QN(n522) );
  DFFX1 \exePacket2_reg[28]  ( .D(n164), .CLK(clk), .Q(computedAddr2_o[27]), 
        .QN(n521) );
  DFFX1 \exePacket2_reg[27]  ( .D(n163), .CLK(clk), .Q(computedAddr2_o[26]), 
        .QN(n520) );
  DFFX1 \exePacket2_reg[26]  ( .D(n162), .CLK(clk), .Q(computedAddr2_o[25]), 
        .QN(n519) );
  DFFX1 \exePacket2_reg[25]  ( .D(n161), .CLK(clk), .Q(computedAddr2_o[24]), 
        .QN(n518) );
  DFFX1 \exePacket2_reg[24]  ( .D(n160), .CLK(clk), .Q(computedAddr2_o[23]), 
        .QN(n517) );
  DFFX1 \exePacket2_reg[23]  ( .D(n159), .CLK(clk), .Q(computedAddr2_o[22]), 
        .QN(n516) );
  DFFX1 \exePacket2_reg[22]  ( .D(n158), .CLK(clk), .Q(computedAddr2_o[21]), 
        .QN(n515) );
  DFFX1 \exePacket2_reg[21]  ( .D(n157), .CLK(clk), .Q(computedAddr2_o[20]), 
        .QN(n514) );
  DFFX1 \exePacket2_reg[20]  ( .D(n156), .CLK(clk), .Q(computedAddr2_o[19]), 
        .QN(n513) );
  DFFX1 \exePacket2_reg[19]  ( .D(n155), .CLK(clk), .Q(computedAddr2_o[18]), 
        .QN(n512) );
  DFFX1 \exePacket2_reg[18]  ( .D(n154), .CLK(clk), .Q(computedAddr2_o[17]), 
        .QN(n511) );
  DFFX1 \exePacket2_reg[17]  ( .D(n153), .CLK(clk), .Q(computedAddr2_o[16]), 
        .QN(n510) );
  DFFX1 \exePacket2_reg[16]  ( .D(n152), .CLK(clk), .Q(computedAddr2_o[15]), 
        .QN(n509) );
  DFFX1 \exePacket2_reg[15]  ( .D(n151), .CLK(clk), .Q(computedAddr2_o[14]), 
        .QN(n508) );
  DFFX1 \exePacket2_reg[14]  ( .D(n150), .CLK(clk), .Q(computedAddr2_o[13]), 
        .QN(n507) );
  DFFX1 \exePacket2_reg[13]  ( .D(n149), .CLK(clk), .Q(computedAddr2_o[12]), 
        .QN(n506) );
  DFFX1 \exePacket2_reg[12]  ( .D(n148), .CLK(clk), .Q(computedAddr2_o[11]), 
        .QN(n505) );
  DFFX1 \exePacket2_reg[11]  ( .D(n147), .CLK(clk), .Q(computedAddr2_o[10]), 
        .QN(n504) );
  DFFX1 \exePacket2_reg[10]  ( .D(n146), .CLK(clk), .Q(computedAddr2_o[9]), 
        .QN(n503) );
  DFFX1 \exePacket2_reg[9]  ( .D(n145), .CLK(clk), .Q(computedAddr2_o[8]), 
        .QN(n502) );
  DFFX1 \exePacket2_reg[8]  ( .D(n144), .CLK(clk), .Q(computedAddr2_o[7]), 
        .QN(n501) );
  DFFX1 \exePacket2_reg[7]  ( .D(n143), .CLK(clk), .Q(computedAddr2_o[6]), 
        .QN(n500) );
  DFFX1 \exePacket2_reg[6]  ( .D(n142), .CLK(clk), .Q(computedAddr2_o[5]), 
        .QN(n499) );
  DFFX1 \exePacket2_reg[5]  ( .D(n141), .CLK(clk), .Q(computedAddr2_o[4]), 
        .QN(n498) );
  DFFX1 \exePacket2_reg[4]  ( .D(n140), .CLK(clk), .Q(computedAddr2_o[3]), 
        .QN(n497) );
  DFFX1 \exePacket2_reg[3]  ( .D(n139), .CLK(clk), .Q(computedAddr2_o[2]), 
        .QN(n496) );
  DFFX1 \exePacket2_reg[2]  ( .D(n138), .CLK(clk), .Q(computedAddr2_o[1]), 
        .QN(n495) );
  DFFX1 \exePacket2_reg[1]  ( .D(n137), .CLK(clk), .Q(computedAddr2_o[0]), 
        .QN(n494) );
  DFFX1 \exePacket2_reg[0]  ( .D(n136), .CLK(clk), .Q(ctrlBrDirection_o) );
  DFFX1 \ldViolationPacket_reg[7]  ( .D(n135), .CLK(clk), .Q(
        ldViolationPacket_o[7]) );
  DFFX1 \ldViolationPacket_reg[6]  ( .D(n134), .CLK(clk), .Q(
        ldViolationPacket_o[6]) );
  DFFX1 \ldViolationPacket_reg[5]  ( .D(n133), .CLK(clk), .Q(
        ldViolationPacket_o[5]) );
  DFFX1 \ldViolationPacket_reg[4]  ( .D(n132), .CLK(clk), .Q(
        ldViolationPacket_o[4]) );
  DFFX1 \ldViolationPacket_reg[3]  ( .D(n131), .CLK(clk), .Q(
        ldViolationPacket_o[3]) );
  DFFX1 \ldViolationPacket_reg[2]  ( .D(n130), .CLK(clk), .Q(
        ldViolationPacket_o[2]) );
  DFFX1 \ldViolationPacket_reg[1]  ( .D(n129), .CLK(clk), .Q(
        ldViolationPacket_o[1]) );
  DFFX1 \ldViolationPacket_reg[0]  ( .D(n128), .CLK(clk), .Q(
        ldViolationPacket_o[0]) );
  DFFX1 \exePacket0_reg[102]  ( .D(n127), .CLK(clk), .Q(ctrlFU0_o[7]) );
  DFFX1 \exePacket0_reg[101]  ( .D(n126), .CLK(clk), .Q(ctrlFU0_o[6]) );
  DFFX1 \exePacket0_reg[100]  ( .D(n125), .CLK(clk), .Q(ctrlFU0_o[5]) );
  DFFX1 \exePacket0_reg[99]  ( .D(n124), .CLK(clk), .Q(ctrlFU0_o[4]) );
  DFFX1 \exePacket0_reg[98]  ( .D(n123), .CLK(clk), .Q(ctrlFU0_o[3]) );
  DFFX1 \exePacket0_reg[97]  ( .D(n122), .CLK(clk), .Q(ctrlFU0_o[2]) );
  DFFX1 \exePacket0_reg[96]  ( .D(n121), .CLK(clk), .Q(ctrlFU0_o[1]) );
  DFFX1 \exePacket0_reg[95]  ( .D(n120), .CLK(clk), .Q(ctrlFU0_o[0]) );
  DFFX1 \exePacket0_reg[94]  ( .D(n119), .CLK(clk), .Q(bypassPacket0_o[41]) );
  DFFX1 \exePacket0_reg[93]  ( .D(n118), .CLK(clk), .Q(bypassPacket0_o[40]) );
  DFFX1 \exePacket0_reg[92]  ( .D(n117), .CLK(clk), .Q(bypassPacket0_o[39]) );
  DFFX1 \exePacket0_reg[91]  ( .D(n116), .CLK(clk), .Q(bypassPacket0_o[38]) );
  DFFX1 \exePacket0_reg[90]  ( .D(n115), .CLK(clk), .Q(bypassPacket0_o[37]) );
  DFFX1 \exePacket0_reg[89]  ( .D(n114), .CLK(clk), .Q(bypassPacket0_o[36]) );
  DFFX1 \exePacket0_reg[88]  ( .D(n113), .CLK(clk), .Q(bypassPacket0_o[35]) );
  DFFX1 \exePacket0_reg[87]  ( .D(n112), .CLK(clk), .Q(ctrlFU0_o[14]) );
  DFFX1 \exePacket0_reg[86]  ( .D(n111), .CLK(clk), .Q(ctrlFU0_o[13]) );
  DFFX1 \exePacket0_reg[85]  ( .D(n110), .CLK(clk), .Q(ctrlFU0_o[12]) );
  DFFX1 \exePacket0_reg[84]  ( .D(n109), .CLK(clk), .Q(ctrlFU0_o[11]) );
  DFFX1 \exePacket0_reg[83]  ( .D(n108), .CLK(clk), .Q(ctrlFU0_o[10]) );
  DFFX1 \exePacket0_reg[82]  ( .D(n107), .CLK(clk), .Q(ctrlFU0_o[9]) );
  DFFX1 \exePacket0_reg[81]  ( .D(n106), .CLK(clk), .Q(ctrlFU0_o[8]) );
  DFFX1 \exePacket0_reg[80]  ( .D(n105), .CLK(clk), .Q(bypassPacket0_o[34]) );
  DFFX1 \exePacket0_reg[79]  ( .D(n104), .CLK(clk), .Q(bypassPacket0_o[33]) );
  DFFX1 \exePacket0_reg[78]  ( .D(n103), .CLK(clk), .Q(bypassPacket0_o[32]) );
  DFFX1 \exePacket0_reg[77]  ( .D(n102), .CLK(clk), .Q(bypassPacket0_o[31]) );
  DFFX1 \exePacket0_reg[76]  ( .D(n101), .CLK(clk), .Q(bypassPacket0_o[30]) );
  DFFX1 \exePacket0_reg[75]  ( .D(n100), .CLK(clk), .Q(bypassPacket0_o[29]) );
  DFFX1 \exePacket0_reg[74]  ( .D(n99), .CLK(clk), .Q(bypassPacket0_o[28]) );
  DFFX1 \exePacket0_reg[73]  ( .D(n98), .CLK(clk), .Q(bypassPacket0_o[27]) );
  DFFX1 \exePacket0_reg[72]  ( .D(n97), .CLK(clk), .Q(bypassPacket0_o[26]) );
  DFFX1 \exePacket0_reg[71]  ( .D(n96), .CLK(clk), .Q(bypassPacket0_o[25]) );
  DFFX1 \exePacket0_reg[70]  ( .D(n95), .CLK(clk), .Q(bypassPacket0_o[24]) );
  DFFX1 \exePacket0_reg[69]  ( .D(n94), .CLK(clk), .Q(bypassPacket0_o[23]) );
  DFFX1 \exePacket0_reg[68]  ( .D(n93), .CLK(clk), .Q(bypassPacket0_o[22]) );
  DFFX1 \exePacket0_reg[67]  ( .D(n92), .CLK(clk), .Q(bypassPacket0_o[21]) );
  DFFX1 \exePacket0_reg[66]  ( .D(n91), .CLK(clk), .Q(bypassPacket0_o[20]) );
  DFFX1 \exePacket0_reg[65]  ( .D(n90), .CLK(clk), .Q(bypassPacket0_o[19]) );
  DFFX1 \exePacket0_reg[64]  ( .D(n89), .CLK(clk), .Q(bypassPacket0_o[18]) );
  DFFX1 \exePacket0_reg[63]  ( .D(n88), .CLK(clk), .Q(bypassPacket0_o[17]) );
  DFFX1 \exePacket0_reg[62]  ( .D(n87), .CLK(clk), .Q(bypassPacket0_o[16]) );
  DFFX1 \exePacket0_reg[61]  ( .D(n86), .CLK(clk), .Q(bypassPacket0_o[15]) );
  DFFX1 \exePacket0_reg[60]  ( .D(n85), .CLK(clk), .Q(bypassPacket0_o[14]) );
  DFFX1 \exePacket0_reg[59]  ( .D(n84), .CLK(clk), .Q(bypassPacket0_o[13]) );
  DFFX1 \exePacket0_reg[58]  ( .D(n83), .CLK(clk), .Q(bypassPacket0_o[12]) );
  DFFX1 \exePacket0_reg[57]  ( .D(n82), .CLK(clk), .Q(bypassPacket0_o[11]) );
  DFFX1 \exePacket0_reg[56]  ( .D(n81), .CLK(clk), .Q(bypassPacket0_o[10]) );
  DFFX1 \exePacket0_reg[55]  ( .D(n80), .CLK(clk), .Q(bypassPacket0_o[9]) );
  DFFX1 \exePacket0_reg[54]  ( .D(n79), .CLK(clk), .Q(bypassPacket0_o[8]) );
  DFFX1 \exePacket0_reg[53]  ( .D(n78), .CLK(clk), .Q(bypassPacket0_o[7]) );
  DFFX1 \exePacket0_reg[52]  ( .D(n77), .CLK(clk), .Q(bypassPacket0_o[6]) );
  DFFX1 \exePacket0_reg[51]  ( .D(n76), .CLK(clk), .Q(bypassPacket0_o[5]) );
  DFFX1 \exePacket0_reg[50]  ( .D(n75), .CLK(clk), .Q(bypassPacket0_o[4]) );
  DFFX1 \exePacket0_reg[49]  ( .D(n74), .CLK(clk), .Q(bypassPacket0_o[3]) );
  DFFX1 \exePacket0_reg[38]  ( .D(n73), .CLK(clk), .Q(bypassPacket0_o[2]) );
  DFFX1 \exePacket0_reg[37]  ( .D(n72), .CLK(clk), .Q(bypassPacket0_o[1]) );
  DFFSSRX1 exePacketValid0_reg ( .D(n6), .RSTB(exePacketValid0_i), .SETB(1'b1), 
        .CLK(clk), .Q(exePacketValid0) );
  DFFX1 \exePacket1_reg[102]  ( .D(n71), .CLK(clk), .Q(ctrlFU1_o[7]) );
  DFFX1 \exePacket1_reg[101]  ( .D(n70), .CLK(clk), .Q(ctrlFU1_o[6]) );
  DFFX1 \exePacket1_reg[100]  ( .D(n69), .CLK(clk), .Q(ctrlFU1_o[5]) );
  DFFX1 \exePacket1_reg[99]  ( .D(n68), .CLK(clk), .Q(ctrlFU1_o[4]) );
  DFFX1 \exePacket1_reg[98]  ( .D(n67), .CLK(clk), .Q(ctrlFU1_o[3]) );
  DFFX1 \exePacket1_reg[97]  ( .D(n66), .CLK(clk), .Q(ctrlFU1_o[2]) );
  DFFX1 \exePacket1_reg[96]  ( .D(n65), .CLK(clk), .Q(ctrlFU1_o[1]) );
  DFFX1 \exePacket1_reg[95]  ( .D(n64), .CLK(clk), .Q(ctrlFU1_o[0]) );
  DFFX1 \exePacket1_reg[94]  ( .D(n63), .CLK(clk), .Q(bypassPacket1_o[41]) );
  DFFX1 \exePacket1_reg[93]  ( .D(n62), .CLK(clk), .Q(bypassPacket1_o[40]) );
  DFFX1 \exePacket1_reg[92]  ( .D(n61), .CLK(clk), .Q(bypassPacket1_o[39]) );
  DFFX1 \exePacket1_reg[91]  ( .D(n60), .CLK(clk), .Q(bypassPacket1_o[38]) );
  DFFX1 \exePacket1_reg[90]  ( .D(n59), .CLK(clk), .Q(bypassPacket1_o[37]) );
  DFFX1 \exePacket1_reg[89]  ( .D(n58), .CLK(clk), .Q(bypassPacket1_o[36]) );
  DFFX1 \exePacket1_reg[88]  ( .D(n57), .CLK(clk), .Q(bypassPacket1_o[35]) );
  DFFX1 \exePacket1_reg[87]  ( .D(n56), .CLK(clk), .Q(ctrlFU1_o[14]) );
  DFFX1 \exePacket1_reg[86]  ( .D(n55), .CLK(clk), .Q(ctrlFU1_o[13]) );
  DFFX1 \exePacket1_reg[85]  ( .D(n54), .CLK(clk), .Q(ctrlFU1_o[12]) );
  DFFX1 \exePacket1_reg[84]  ( .D(n53), .CLK(clk), .Q(ctrlFU1_o[11]) );
  DFFX1 \exePacket1_reg[83]  ( .D(n52), .CLK(clk), .Q(ctrlFU1_o[10]) );
  DFFX1 \exePacket1_reg[82]  ( .D(n51), .CLK(clk), .Q(ctrlFU1_o[9]) );
  DFFX1 \exePacket1_reg[81]  ( .D(n50), .CLK(clk), .Q(ctrlFU1_o[8]) );
  DFFX1 \exePacket1_reg[80]  ( .D(n49), .CLK(clk), .Q(bypassPacket1_o[34]) );
  DFFX1 \exePacket1_reg[79]  ( .D(n48), .CLK(clk), .Q(bypassPacket1_o[33]) );
  DFFX1 \exePacket1_reg[78]  ( .D(n47), .CLK(clk), .Q(bypassPacket1_o[32]) );
  DFFX1 \exePacket1_reg[77]  ( .D(n46), .CLK(clk), .Q(bypassPacket1_o[31]) );
  DFFX1 \exePacket1_reg[76]  ( .D(n45), .CLK(clk), .Q(bypassPacket1_o[30]) );
  DFFX1 \exePacket1_reg[75]  ( .D(n44), .CLK(clk), .Q(bypassPacket1_o[29]) );
  DFFX1 \exePacket1_reg[74]  ( .D(n43), .CLK(clk), .Q(bypassPacket1_o[28]) );
  DFFX1 \exePacket1_reg[73]  ( .D(n42), .CLK(clk), .Q(bypassPacket1_o[27]) );
  DFFX1 \exePacket1_reg[72]  ( .D(n41), .CLK(clk), .Q(bypassPacket1_o[26]) );
  DFFX1 \exePacket1_reg[71]  ( .D(n40), .CLK(clk), .Q(bypassPacket1_o[25]) );
  DFFX1 \exePacket1_reg[70]  ( .D(n39), .CLK(clk), .Q(bypassPacket1_o[24]) );
  DFFX1 \exePacket1_reg[69]  ( .D(n38), .CLK(clk), .Q(bypassPacket1_o[23]) );
  DFFX1 \exePacket1_reg[68]  ( .D(n37), .CLK(clk), .Q(bypassPacket1_o[22]) );
  DFFX1 \exePacket1_reg[67]  ( .D(n36), .CLK(clk), .Q(bypassPacket1_o[21]) );
  DFFX1 \exePacket1_reg[66]  ( .D(n35), .CLK(clk), .Q(bypassPacket1_o[20]) );
  DFFX1 \exePacket1_reg[65]  ( .D(n34), .CLK(clk), .Q(bypassPacket1_o[19]) );
  DFFX1 \exePacket1_reg[64]  ( .D(n33), .CLK(clk), .Q(bypassPacket1_o[18]) );
  DFFX1 \exePacket1_reg[63]  ( .D(n32), .CLK(clk), .Q(bypassPacket1_o[17]) );
  DFFX1 \exePacket1_reg[62]  ( .D(n31), .CLK(clk), .Q(bypassPacket1_o[16]) );
  DFFX1 \exePacket1_reg[61]  ( .D(n30), .CLK(clk), .Q(bypassPacket1_o[15]) );
  DFFX1 \exePacket1_reg[60]  ( .D(n29), .CLK(clk), .Q(bypassPacket1_o[14]) );
  DFFX1 \exePacket1_reg[59]  ( .D(n28), .CLK(clk), .Q(bypassPacket1_o[13]) );
  DFFX1 \exePacket1_reg[58]  ( .D(n27), .CLK(clk), .Q(bypassPacket1_o[12]) );
  DFFX1 \exePacket1_reg[57]  ( .D(n26), .CLK(clk), .Q(bypassPacket1_o[11]) );
  DFFX1 \exePacket1_reg[56]  ( .D(n25), .CLK(clk), .Q(bypassPacket1_o[10]) );
  DFFX1 \exePacket1_reg[55]  ( .D(n24), .CLK(clk), .Q(bypassPacket1_o[9]) );
  DFFX1 \exePacket1_reg[54]  ( .D(n23), .CLK(clk), .Q(bypassPacket1_o[8]) );
  DFFX1 \exePacket1_reg[53]  ( .D(n22), .CLK(clk), .Q(bypassPacket1_o[7]) );
  DFFX1 \exePacket1_reg[52]  ( .D(n21), .CLK(clk), .Q(bypassPacket1_o[6]) );
  DFFX1 \exePacket1_reg[51]  ( .D(n20), .CLK(clk), .Q(bypassPacket1_o[5]) );
  DFFX1 \exePacket1_reg[50]  ( .D(n19), .CLK(clk), .Q(bypassPacket1_o[4]) );
  DFFX1 \exePacket1_reg[49]  ( .D(n18), .CLK(clk), .Q(bypassPacket1_o[3]) );
  DFFX1 \exePacket1_reg[38]  ( .D(n17), .CLK(clk), .Q(bypassPacket1_o[2]) );
  DFFX1 \exePacket1_reg[37]  ( .D(n16), .CLK(clk), .Q(bypassPacket1_o[1]) );
  AO22X1 U18 ( .IN1(bypassPacket2_o[29]), .IN2(n593), .IN3(exePacket2_i[75]), 
        .IN4(n584), .Q(n201) );
  AO22X1 U19 ( .IN1(bypassPacket2_o[30]), .IN2(n593), .IN3(exePacket2_i[76]), 
        .IN4(n8), .Q(n202) );
  AO22X1 U20 ( .IN1(bypassPacket2_o[31]), .IN2(n593), .IN3(exePacket2_i[77]), 
        .IN4(n8), .Q(n203) );
  AO22X1 U21 ( .IN1(bypassPacket2_o[32]), .IN2(n593), .IN3(exePacket2_i[78]), 
        .IN4(n585), .Q(n204) );
  AO22X1 U22 ( .IN1(bypassPacket2_o[33]), .IN2(n593), .IN3(exePacket2_i[79]), 
        .IN4(n587), .Q(n205) );
  AO22X1 U23 ( .IN1(bypassPacket2_o[34]), .IN2(n593), .IN3(exePacket2_i[80]), 
        .IN4(n586), .Q(n206) );
  AO22X1 U24 ( .IN1(ctrlFU2_o[8]), .IN2(n593), .IN3(exePacket2_i[81]), .IN4(
        n587), .Q(n207) );
  AO22X1 U25 ( .IN1(ctrlFU2_o[9]), .IN2(n593), .IN3(exePacket2_i[82]), .IN4(
        n586), .Q(n208) );
  AO22X1 U26 ( .IN1(ctrlFU2_o[10]), .IN2(n593), .IN3(exePacket2_i[83]), .IN4(
        n585), .Q(n209) );
  AO22X1 U27 ( .IN1(ctrlFU2_o[11]), .IN2(n593), .IN3(exePacket2_i[84]), .IN4(
        n585), .Q(n210) );
  AO22X1 U28 ( .IN1(ctrlFU2_o[12]), .IN2(n589), .IN3(exePacket2_i[85]), .IN4(
        n584), .Q(n211) );
  AO22X1 U29 ( .IN1(ctrlFU2_o[13]), .IN2(n588), .IN3(exePacket2_i[86]), .IN4(
        n8), .Q(n212) );
  AO22X1 U30 ( .IN1(ctrlFU2_o[14]), .IN2(n590), .IN3(exePacket2_i[87]), .IN4(
        n8), .Q(n213) );
  AO22X1 U31 ( .IN1(bypassPacket2_o[35]), .IN2(n591), .IN3(exePacket2_i[88]), 
        .IN4(n587), .Q(n214) );
  AO22X1 U32 ( .IN1(bypassPacket2_o[36]), .IN2(n592), .IN3(exePacket2_i[89]), 
        .IN4(n586), .Q(n215) );
  AO22X1 U33 ( .IN1(bypassPacket2_o[37]), .IN2(n588), .IN3(exePacket2_i[90]), 
        .IN4(n585), .Q(n216) );
  AO22X1 U34 ( .IN1(bypassPacket2_o[38]), .IN2(n593), .IN3(exePacket2_i[91]), 
        .IN4(n584), .Q(n217) );
  AO22X1 U35 ( .IN1(bypassPacket2_o[39]), .IN2(n589), .IN3(exePacket2_i[92]), 
        .IN4(n8), .Q(n218) );
  AO22X1 U36 ( .IN1(bypassPacket2_o[40]), .IN2(n588), .IN3(exePacket2_i[93]), 
        .IN4(n8), .Q(n219) );
  AO22X1 U37 ( .IN1(bypassPacket2_o[41]), .IN2(n590), .IN3(exePacket2_i[94]), 
        .IN4(n587), .Q(n220) );
  AO22X1 U38 ( .IN1(ctrlFU2_o[0]), .IN2(n591), .IN3(exePacket2_i[95]), .IN4(
        n586), .Q(n221) );
  AO22X1 U39 ( .IN1(ctrlFU2_o[1]), .IN2(n592), .IN3(exePacket2_i[96]), .IN4(
        n584), .Q(n222) );
  AO22X1 U40 ( .IN1(ctrlFU2_o[2]), .IN2(n589), .IN3(exePacket2_i[97]), .IN4(n8), .Q(n223) );
  AO22X1 U41 ( .IN1(ctrlFU2_o[3]), .IN2(n593), .IN3(exePacket2_i[98]), .IN4(
        n587), .Q(n224) );
  AO22X1 U42 ( .IN1(ctrlFU2_o[4]), .IN2(n589), .IN3(exePacket2_i[99]), .IN4(
        n586), .Q(n225) );
  AO22X1 U43 ( .IN1(ctrlFU2_o[5]), .IN2(n588), .IN3(exePacket2_i[100]), .IN4(
        n585), .Q(n226) );
  AO22X1 U44 ( .IN1(ctrlFU2_o[6]), .IN2(n593), .IN3(exePacket2_i[101]), .IN4(
        n584), .Q(n227) );
  AO22X1 U45 ( .IN1(ctrlFU2_o[7]), .IN2(n590), .IN3(exePacket2_i[102]), .IN4(
        n8), .Q(n228) );
  AO22X1 U46 ( .IN1(agenIqEntry0_o[0]), .IN2(n583), .IN3(lsuPacket0_i[0]), 
        .IN4(n10), .Q(n229) );
  AO22X1 U47 ( .IN1(agenIqEntry0_o[1]), .IN2(n583), .IN3(lsuPacket0_i[1]), 
        .IN4(n10), .Q(n230) );
  AO22X1 U48 ( .IN1(agenIqEntry0_o[2]), .IN2(n583), .IN3(lsuPacket0_i[2]), 
        .IN4(n10), .Q(n231) );
  AO22X1 U49 ( .IN1(agenIqEntry0_o[3]), .IN2(n583), .IN3(lsuPacket0_i[3]), 
        .IN4(n10), .Q(n232) );
  AO22X1 U50 ( .IN1(agenIqEntry0_o[4]), .IN2(n583), .IN3(lsuPacket0_i[4]), 
        .IN4(n10), .Q(n233) );
  AO22X1 U51 ( .IN1(ctrlFU3_o[8]), .IN2(n583), .IN3(lsuPacket0_i[5]), .IN4(n10), .Q(n234) );
  AO22X1 U52 ( .IN1(ctrlFU3_o[9]), .IN2(n583), .IN3(lsuPacket0_i[6]), .IN4(
        n581), .Q(n235) );
  AO22X1 U53 ( .IN1(ctrlFU3_o[10]), .IN2(n583), .IN3(lsuPacket0_i[7]), .IN4(
        n580), .Q(n236) );
  AO22X1 U54 ( .IN1(ctrlFU3_o[11]), .IN2(n583), .IN3(lsuPacket0_i[8]), .IN4(
        n579), .Q(n237) );
  AO22X1 U55 ( .IN1(ctrlFU3_o[12]), .IN2(n583), .IN3(lsuPacket0_i[9]), .IN4(
        n581), .Q(n238) );
  AO22X1 U56 ( .IN1(ctrlFU3_o[13]), .IN2(n583), .IN3(lsuPacket0_i[10]), .IN4(
        n580), .Q(n239) );
  AO22X1 U57 ( .IN1(ctrlFU3_o[14]), .IN2(n583), .IN3(lsuPacket0_i[11]), .IN4(
        n579), .Q(n240) );
  AO22X1 U58 ( .IN1(bypassPacket3_o[35]), .IN2(n9), .IN3(lsuPacket0_i[12]), 
        .IN4(n10), .Q(n241) );
  AO22X1 U59 ( .IN1(bypassPacket3_o[36]), .IN2(n583), .IN3(lsuPacket0_i[13]), 
        .IN4(n10), .Q(n242) );
  AO22X1 U60 ( .IN1(bypassPacket3_o[37]), .IN2(n9), .IN3(lsuPacket0_i[14]), 
        .IN4(n10), .Q(n243) );
  AO22X1 U61 ( .IN1(bypassPacket3_o[38]), .IN2(n583), .IN3(lsuPacket0_i[15]), 
        .IN4(n581), .Q(n244) );
  AO22X1 U62 ( .IN1(bypassPacket3_o[39]), .IN2(n583), .IN3(lsuPacket0_i[16]), 
        .IN4(n580), .Q(n245) );
  AO22X1 U63 ( .IN1(bypassPacket3_o[40]), .IN2(n583), .IN3(lsuPacket0_i[17]), 
        .IN4(n579), .Q(n246) );
  AO22X1 U64 ( .IN1(bypassPacket3_o[41]), .IN2(n583), .IN3(lsuPacket0_i[18]), 
        .IN4(n10), .Q(n247) );
  AO22X1 U65 ( .IN1(bypassPacket3_o[3]), .IN2(n583), .IN3(lsuPacket0_i[19]), 
        .IN4(n581), .Q(n248) );
  AO22X1 U66 ( .IN1(bypassPacket3_o[4]), .IN2(n583), .IN3(lsuPacket0_i[20]), 
        .IN4(n580), .Q(n249) );
  AO22X1 U67 ( .IN1(bypassPacket3_o[5]), .IN2(n583), .IN3(lsuPacket0_i[21]), 
        .IN4(n579), .Q(n250) );
  AO22X1 U68 ( .IN1(bypassPacket3_o[6]), .IN2(n9), .IN3(lsuPacket0_i[22]), 
        .IN4(n10), .Q(n251) );
  AO22X1 U69 ( .IN1(bypassPacket3_o[7]), .IN2(n583), .IN3(lsuPacket0_i[23]), 
        .IN4(n581), .Q(n252) );
  AO22X1 U70 ( .IN1(bypassPacket3_o[8]), .IN2(n9), .IN3(lsuPacket0_i[24]), 
        .IN4(n579), .Q(n253) );
  AO22X1 U71 ( .IN1(bypassPacket3_o[9]), .IN2(n9), .IN3(lsuPacket0_i[25]), 
        .IN4(n579), .Q(n254) );
  AO22X1 U72 ( .IN1(bypassPacket3_o[10]), .IN2(n9), .IN3(lsuPacket0_i[26]), 
        .IN4(n579), .Q(n255) );
  AO22X1 U73 ( .IN1(bypassPacket3_o[11]), .IN2(n9), .IN3(lsuPacket0_i[27]), 
        .IN4(n579), .Q(n256) );
  AO22X1 U74 ( .IN1(bypassPacket3_o[12]), .IN2(n582), .IN3(lsuPacket0_i[28]), 
        .IN4(n579), .Q(n257) );
  AO22X1 U75 ( .IN1(bypassPacket3_o[13]), .IN2(n583), .IN3(lsuPacket0_i[29]), 
        .IN4(n579), .Q(n258) );
  AO22X1 U76 ( .IN1(bypassPacket3_o[14]), .IN2(n583), .IN3(lsuPacket0_i[30]), 
        .IN4(n579), .Q(n259) );
  AO22X1 U77 ( .IN1(bypassPacket3_o[15]), .IN2(n583), .IN3(lsuPacket0_i[31]), 
        .IN4(n579), .Q(n260) );
  AO22X1 U78 ( .IN1(bypassPacket3_o[16]), .IN2(n583), .IN3(lsuPacket0_i[32]), 
        .IN4(n579), .Q(n261) );
  AO22X1 U79 ( .IN1(bypassPacket3_o[17]), .IN2(n583), .IN3(lsuPacket0_i[33]), 
        .IN4(n579), .Q(n262) );
  AO22X1 U80 ( .IN1(bypassPacket3_o[18]), .IN2(n583), .IN3(lsuPacket0_i[34]), 
        .IN4(n579), .Q(n263) );
  AO22X1 U81 ( .IN1(bypassPacket3_o[19]), .IN2(n583), .IN3(lsuPacket0_i[35]), 
        .IN4(n579), .Q(n264) );
  AO22X1 U82 ( .IN1(bypassPacket3_o[20]), .IN2(n9), .IN3(lsuPacket0_i[36]), 
        .IN4(n580), .Q(n265) );
  AO22X1 U83 ( .IN1(bypassPacket3_o[21]), .IN2(n9), .IN3(lsuPacket0_i[37]), 
        .IN4(n580), .Q(n266) );
  AO22X1 U84 ( .IN1(bypassPacket3_o[22]), .IN2(n9), .IN3(lsuPacket0_i[38]), 
        .IN4(n580), .Q(n267) );
  AO22X1 U85 ( .IN1(bypassPacket3_o[23]), .IN2(n9), .IN3(lsuPacket0_i[39]), 
        .IN4(n580), .Q(n268) );
  AO22X1 U86 ( .IN1(bypassPacket3_o[24]), .IN2(n9), .IN3(lsuPacket0_i[40]), 
        .IN4(n580), .Q(n269) );
  AO22X1 U87 ( .IN1(bypassPacket3_o[25]), .IN2(n9), .IN3(lsuPacket0_i[41]), 
        .IN4(n580), .Q(n270) );
  AO22X1 U88 ( .IN1(bypassPacket3_o[26]), .IN2(n9), .IN3(lsuPacket0_i[42]), 
        .IN4(n580), .Q(n271) );
  AO22X1 U89 ( .IN1(bypassPacket3_o[27]), .IN2(n582), .IN3(lsuPacket0_i[43]), 
        .IN4(n580), .Q(n272) );
  AO22X1 U90 ( .IN1(bypassPacket3_o[28]), .IN2(n582), .IN3(lsuPacket0_i[44]), 
        .IN4(n580), .Q(n273) );
  AO22X1 U91 ( .IN1(bypassPacket3_o[29]), .IN2(n582), .IN3(lsuPacket0_i[45]), 
        .IN4(n580), .Q(n274) );
  AO22X1 U92 ( .IN1(bypassPacket3_o[30]), .IN2(n582), .IN3(lsuPacket0_i[46]), 
        .IN4(n580), .Q(n275) );
  AO22X1 U93 ( .IN1(bypassPacket3_o[31]), .IN2(n582), .IN3(lsuPacket0_i[47]), 
        .IN4(n580), .Q(n276) );
  AO22X1 U94 ( .IN1(bypassPacket3_o[32]), .IN2(n582), .IN3(lsuPacket0_i[48]), 
        .IN4(n581), .Q(n277) );
  AO22X1 U95 ( .IN1(bypassPacket3_o[33]), .IN2(n582), .IN3(lsuPacket0_i[49]), 
        .IN4(n581), .Q(n278) );
  AO22X1 U96 ( .IN1(bypassPacket3_o[34]), .IN2(n582), .IN3(lsuPacket0_i[50]), 
        .IN4(n581), .Q(n279) );
  AO22X1 U97 ( .IN1(ctrlFU3_o[0]), .IN2(n582), .IN3(lsuPacket0_i[51]), .IN4(
        n581), .Q(n280) );
  AO22X1 U98 ( .IN1(ctrlFU3_o[1]), .IN2(n582), .IN3(lsuPacket0_i[52]), .IN4(
        n581), .Q(n281) );
  AO22X1 U99 ( .IN1(ctrlFU3_o[2]), .IN2(n582), .IN3(lsuPacket0_i[53]), .IN4(
        n581), .Q(n282) );
  AO22X1 U100 ( .IN1(ctrlFU3_o[3]), .IN2(n582), .IN3(lsuPacket0_i[54]), .IN4(
        n581), .Q(n283) );
  AO22X1 U101 ( .IN1(ctrlFU3_o[4]), .IN2(n582), .IN3(lsuPacket0_i[55]), .IN4(
        n581), .Q(n284) );
  AO22X1 U102 ( .IN1(ctrlFU3_o[5]), .IN2(n582), .IN3(lsuPacket0_i[56]), .IN4(
        n581), .Q(n285) );
  AO22X1 U103 ( .IN1(ctrlFU3_o[6]), .IN2(n582), .IN3(lsuPacket0_i[57]), .IN4(
        n581), .Q(n286) );
  AO22X1 U104 ( .IN1(ctrlFU3_o[7]), .IN2(n582), .IN3(lsuPacket0_i[58]), .IN4(
        n581), .Q(n287) );
  AO22X1 U105 ( .IN1(bypassPacket1_o[1]), .IN2(n578), .IN3(exePacket1_i_37), 
        .IN4(n574), .Q(n16) );
  AO22X1 U106 ( .IN1(bypassPacket1_o[2]), .IN2(n578), .IN3(exePacket1_i_38), 
        .IN4(n574), .Q(n17) );
  AO22X1 U107 ( .IN1(bypassPacket1_o[3]), .IN2(n578), .IN3(exePacket1_i[49]), 
        .IN4(n574), .Q(n18) );
  AO22X1 U108 ( .IN1(bypassPacket1_o[4]), .IN2(n578), .IN3(exePacket1_i[50]), 
        .IN4(n574), .Q(n19) );
  AO22X1 U109 ( .IN1(bypassPacket1_o[5]), .IN2(n578), .IN3(exePacket1_i[51]), 
        .IN4(n574), .Q(n20) );
  AO22X1 U110 ( .IN1(bypassPacket1_o[6]), .IN2(n578), .IN3(exePacket1_i[52]), 
        .IN4(n574), .Q(n21) );
  AO22X1 U111 ( .IN1(bypassPacket1_o[7]), .IN2(n578), .IN3(exePacket1_i[53]), 
        .IN4(n574), .Q(n22) );
  AO22X1 U112 ( .IN1(bypassPacket1_o[8]), .IN2(n578), .IN3(exePacket1_i[54]), 
        .IN4(n574), .Q(n23) );
  AO22X1 U113 ( .IN1(bypassPacket1_o[9]), .IN2(n578), .IN3(exePacket1_i[55]), 
        .IN4(n574), .Q(n24) );
  AO22X1 U114 ( .IN1(bypassPacket1_o[10]), .IN2(n578), .IN3(exePacket1_i[56]), 
        .IN4(n574), .Q(n25) );
  AO22X1 U115 ( .IN1(bypassPacket1_o[11]), .IN2(n578), .IN3(exePacket1_i[57]), 
        .IN4(n574), .Q(n26) );
  AO22X1 U116 ( .IN1(bypassPacket1_o[12]), .IN2(n578), .IN3(exePacket1_i[58]), 
        .IN4(n574), .Q(n27) );
  AO22X1 U117 ( .IN1(bypassPacket1_o[13]), .IN2(n578), .IN3(exePacket1_i[59]), 
        .IN4(n575), .Q(n28) );
  AO22X1 U118 ( .IN1(bypassPacket1_o[14]), .IN2(n578), .IN3(exePacket1_i[60]), 
        .IN4(n575), .Q(n29) );
  AO22X1 U119 ( .IN1(bypassPacket1_o[15]), .IN2(n578), .IN3(exePacket1_i[61]), 
        .IN4(n575), .Q(n30) );
  AO22X1 U120 ( .IN1(bypassPacket1_o[16]), .IN2(n578), .IN3(exePacket1_i[62]), 
        .IN4(n575), .Q(n31) );
  AO22X1 U121 ( .IN1(bypassPacket1_o[17]), .IN2(n578), .IN3(exePacket1_i[63]), 
        .IN4(n575), .Q(n32) );
  AO22X1 U122 ( .IN1(bypassPacket1_o[18]), .IN2(n578), .IN3(exePacket1_i[64]), 
        .IN4(n575), .Q(n33) );
  AO22X1 U123 ( .IN1(bypassPacket1_o[19]), .IN2(n578), .IN3(exePacket1_i[65]), 
        .IN4(n575), .Q(n34) );
  AO22X1 U124 ( .IN1(bypassPacket1_o[20]), .IN2(n11), .IN3(exePacket1_i[66]), 
        .IN4(n575), .Q(n35) );
  AO22X1 U125 ( .IN1(bypassPacket1_o[21]), .IN2(n578), .IN3(exePacket1_i[67]), 
        .IN4(n575), .Q(n36) );
  AO22X1 U126 ( .IN1(bypassPacket1_o[22]), .IN2(n578), .IN3(exePacket1_i[68]), 
        .IN4(n575), .Q(n37) );
  AO22X1 U127 ( .IN1(bypassPacket1_o[23]), .IN2(n578), .IN3(exePacket1_i[69]), 
        .IN4(n575), .Q(n38) );
  AO22X1 U128 ( .IN1(bypassPacket1_o[24]), .IN2(n578), .IN3(exePacket1_i[70]), 
        .IN4(n575), .Q(n39) );
  AO22X1 U129 ( .IN1(bypassPacket1_o[25]), .IN2(n11), .IN3(exePacket1_i[71]), 
        .IN4(n12), .Q(n40) );
  AO22X1 U130 ( .IN1(bypassPacket1_o[26]), .IN2(n11), .IN3(exePacket1_i[72]), 
        .IN4(n12), .Q(n41) );
  AO22X1 U131 ( .IN1(bypassPacket1_o[27]), .IN2(n11), .IN3(exePacket1_i[73]), 
        .IN4(n12), .Q(n42) );
  AO22X1 U132 ( .IN1(bypassPacket1_o[28]), .IN2(n11), .IN3(exePacket1_i[74]), 
        .IN4(n12), .Q(n43) );
  AO22X1 U133 ( .IN1(bypassPacket1_o[29]), .IN2(n11), .IN3(exePacket1_i[75]), 
        .IN4(n12), .Q(n44) );
  AO22X1 U134 ( .IN1(bypassPacket1_o[30]), .IN2(n11), .IN3(exePacket1_i[76]), 
        .IN4(n12), .Q(n45) );
  AO22X1 U135 ( .IN1(bypassPacket1_o[31]), .IN2(n578), .IN3(exePacket1_i[77]), 
        .IN4(n575), .Q(n46) );
  AO22X1 U136 ( .IN1(bypassPacket1_o[32]), .IN2(n578), .IN3(exePacket1_i[78]), 
        .IN4(n574), .Q(n47) );
  AO22X1 U137 ( .IN1(bypassPacket1_o[33]), .IN2(n578), .IN3(exePacket1_i[79]), 
        .IN4(n576), .Q(n48) );
  AO22X1 U138 ( .IN1(bypassPacket1_o[34]), .IN2(n578), .IN3(exePacket1_i[80]), 
        .IN4(n575), .Q(n49) );
  AO22X1 U139 ( .IN1(ctrlFU1_o[8]), .IN2(n578), .IN3(exePacket1_i[81]), .IN4(
        n574), .Q(n50) );
  AO22X1 U140 ( .IN1(ctrlFU1_o[9]), .IN2(n577), .IN3(exePacket1_i[82]), .IN4(
        n576), .Q(n51) );
  AO22X1 U141 ( .IN1(ctrlFU1_o[10]), .IN2(n11), .IN3(exePacket1_i[83]), .IN4(
        n576), .Q(n52) );
  AO22X1 U142 ( .IN1(ctrlFU1_o[11]), .IN2(n11), .IN3(exePacket1_i[84]), .IN4(
        n576), .Q(n53) );
  AO22X1 U143 ( .IN1(ctrlFU1_o[12]), .IN2(n11), .IN3(exePacket1_i[85]), .IN4(
        n576), .Q(n54) );
  AO22X1 U144 ( .IN1(ctrlFU1_o[13]), .IN2(n11), .IN3(exePacket1_i[86]), .IN4(
        n576), .Q(n55) );
  AO22X1 U145 ( .IN1(ctrlFU1_o[14]), .IN2(n577), .IN3(exePacket1_i[87]), .IN4(
        n576), .Q(n56) );
  AO22X1 U146 ( .IN1(bypassPacket1_o[35]), .IN2(n577), .IN3(exePacket1_i[88]), 
        .IN4(n12), .Q(n57) );
  AO22X1 U147 ( .IN1(bypassPacket1_o[36]), .IN2(n577), .IN3(exePacket1_i[89]), 
        .IN4(n575), .Q(n58) );
  AO22X1 U148 ( .IN1(bypassPacket1_o[37]), .IN2(n577), .IN3(exePacket1_i[90]), 
        .IN4(n574), .Q(n59) );
  AO22X1 U149 ( .IN1(bypassPacket1_o[38]), .IN2(n577), .IN3(exePacket1_i[91]), 
        .IN4(n576), .Q(n60) );
  AO22X1 U150 ( .IN1(bypassPacket1_o[39]), .IN2(n577), .IN3(exePacket1_i[92]), 
        .IN4(n12), .Q(n61) );
  AO22X1 U151 ( .IN1(bypassPacket1_o[40]), .IN2(n577), .IN3(exePacket1_i[93]), 
        .IN4(n575), .Q(n62) );
  AO22X1 U152 ( .IN1(bypassPacket1_o[41]), .IN2(n577), .IN3(exePacket1_i[94]), 
        .IN4(n574), .Q(n63) );
  AO22X1 U153 ( .IN1(ctrlFU1_o[0]), .IN2(n577), .IN3(exePacket1_i[95]), .IN4(
        n576), .Q(n64) );
  AO22X1 U154 ( .IN1(ctrlFU1_o[1]), .IN2(n577), .IN3(exePacket1_i[96]), .IN4(
        n576), .Q(n65) );
  AO22X1 U155 ( .IN1(ctrlFU1_o[2]), .IN2(n577), .IN3(exePacket1_i[97]), .IN4(
        n576), .Q(n66) );
  AO22X1 U156 ( .IN1(ctrlFU1_o[3]), .IN2(n577), .IN3(exePacket1_i[98]), .IN4(
        n576), .Q(n67) );
  AO22X1 U157 ( .IN1(ctrlFU1_o[4]), .IN2(n577), .IN3(exePacket1_i[99]), .IN4(
        n576), .Q(n68) );
  AO22X1 U158 ( .IN1(ctrlFU1_o[5]), .IN2(n577), .IN3(exePacket1_i[100]), .IN4(
        n576), .Q(n69) );
  AO22X1 U159 ( .IN1(ctrlFU1_o[6]), .IN2(n577), .IN3(exePacket1_i[101]), .IN4(
        n576), .Q(n70) );
  AO22X1 U160 ( .IN1(ctrlFU1_o[7]), .IN2(n577), .IN3(exePacket1_i[102]), .IN4(
        n576), .Q(n71) );
  AO22X1 U161 ( .IN1(bypassPacket0_o[1]), .IN2(n573), .IN3(exePacket0_i_37), 
        .IN4(n570), .Q(n72) );
  AO22X1 U162 ( .IN1(bypassPacket0_o[2]), .IN2(n573), .IN3(exePacket0_i_38), 
        .IN4(n569), .Q(n73) );
  AO22X1 U163 ( .IN1(bypassPacket0_o[3]), .IN2(n572), .IN3(exePacket0_i[49]), 
        .IN4(n568), .Q(n74) );
  AO22X1 U164 ( .IN1(bypassPacket0_o[4]), .IN2(n572), .IN3(exePacket0_i[50]), 
        .IN4(n570), .Q(n75) );
  AO22X1 U165 ( .IN1(bypassPacket0_o[5]), .IN2(n572), .IN3(exePacket0_i[51]), 
        .IN4(n570), .Q(n76) );
  AO22X1 U166 ( .IN1(bypassPacket0_o[6]), .IN2(n572), .IN3(exePacket0_i[52]), 
        .IN4(n569), .Q(n77) );
  AO22X1 U167 ( .IN1(bypassPacket0_o[7]), .IN2(n572), .IN3(exePacket0_i[53]), 
        .IN4(n568), .Q(n78) );
  AO22X1 U168 ( .IN1(bypassPacket0_o[8]), .IN2(n572), .IN3(exePacket0_i[54]), 
        .IN4(n569), .Q(n79) );
  AO22X1 U169 ( .IN1(bypassPacket0_o[9]), .IN2(n572), .IN3(exePacket0_i[55]), 
        .IN4(n568), .Q(n80) );
  AO22X1 U170 ( .IN1(bypassPacket0_o[10]), .IN2(n572), .IN3(exePacket0_i[56]), 
        .IN4(n570), .Q(n81) );
  AO22X1 U171 ( .IN1(bypassPacket0_o[11]), .IN2(n572), .IN3(exePacket0_i[57]), 
        .IN4(n569), .Q(n82) );
  AO22X1 U172 ( .IN1(bypassPacket0_o[12]), .IN2(n572), .IN3(exePacket0_i[58]), 
        .IN4(n568), .Q(n83) );
  AO22X1 U173 ( .IN1(bypassPacket0_o[13]), .IN2(n572), .IN3(exePacket0_i[59]), 
        .IN4(n568), .Q(n84) );
  AO22X1 U174 ( .IN1(bypassPacket0_o[14]), .IN2(n572), .IN3(exePacket0_i[60]), 
        .IN4(n568), .Q(n85) );
  AO22X1 U175 ( .IN1(bypassPacket0_o[15]), .IN2(n572), .IN3(exePacket0_i[61]), 
        .IN4(n568), .Q(n86) );
  AO22X1 U176 ( .IN1(bypassPacket0_o[16]), .IN2(n572), .IN3(exePacket0_i[62]), 
        .IN4(n568), .Q(n87) );
  AO22X1 U177 ( .IN1(bypassPacket0_o[17]), .IN2(n572), .IN3(exePacket0_i[63]), 
        .IN4(n568), .Q(n88) );
  AO22X1 U178 ( .IN1(bypassPacket0_o[18]), .IN2(n572), .IN3(exePacket0_i[64]), 
        .IN4(n568), .Q(n89) );
  AO22X1 U179 ( .IN1(bypassPacket0_o[19]), .IN2(n572), .IN3(exePacket0_i[65]), 
        .IN4(n568), .Q(n90) );
  AO22X1 U180 ( .IN1(bypassPacket0_o[20]), .IN2(n572), .IN3(exePacket0_i[66]), 
        .IN4(n568), .Q(n91) );
  AO22X1 U181 ( .IN1(bypassPacket0_o[21]), .IN2(n572), .IN3(exePacket0_i[67]), 
        .IN4(n568), .Q(n92) );
  AO22X1 U182 ( .IN1(bypassPacket0_o[22]), .IN2(n571), .IN3(exePacket0_i[68]), 
        .IN4(n568), .Q(n93) );
  AO22X1 U183 ( .IN1(bypassPacket0_o[23]), .IN2(n571), .IN3(exePacket0_i[69]), 
        .IN4(n568), .Q(n94) );
  AO22X1 U184 ( .IN1(bypassPacket0_o[24]), .IN2(n571), .IN3(exePacket0_i[70]), 
        .IN4(n568), .Q(n95) );
  AO22X1 U185 ( .IN1(bypassPacket0_o[25]), .IN2(n571), .IN3(exePacket0_i[71]), 
        .IN4(n569), .Q(n96) );
  AO22X1 U186 ( .IN1(bypassPacket0_o[26]), .IN2(n571), .IN3(exePacket0_i[72]), 
        .IN4(n569), .Q(n97) );
  AO22X1 U187 ( .IN1(bypassPacket0_o[27]), .IN2(n571), .IN3(exePacket0_i[73]), 
        .IN4(n569), .Q(n98) );
  AO22X1 U188 ( .IN1(bypassPacket0_o[28]), .IN2(n571), .IN3(exePacket0_i[74]), 
        .IN4(n569), .Q(n99) );
  AO22X1 U189 ( .IN1(bypassPacket0_o[29]), .IN2(n571), .IN3(exePacket0_i[75]), 
        .IN4(n569), .Q(n100) );
  AO22X1 U190 ( .IN1(bypassPacket0_o[30]), .IN2(n571), .IN3(exePacket0_i[76]), 
        .IN4(n569), .Q(n101) );
  AO22X1 U191 ( .IN1(bypassPacket0_o[31]), .IN2(n571), .IN3(exePacket0_i[77]), 
        .IN4(n569), .Q(n102) );
  AO22X1 U192 ( .IN1(bypassPacket0_o[32]), .IN2(n571), .IN3(exePacket0_i[78]), 
        .IN4(n569), .Q(n103) );
  AO22X1 U193 ( .IN1(bypassPacket0_o[33]), .IN2(n571), .IN3(exePacket0_i[79]), 
        .IN4(n569), .Q(n104) );
  AO22X1 U194 ( .IN1(bypassPacket0_o[34]), .IN2(n571), .IN3(exePacket0_i[80]), 
        .IN4(n569), .Q(n105) );
  AO22X1 U195 ( .IN1(ctrlFU0_o[8]), .IN2(n571), .IN3(exePacket0_i[81]), .IN4(
        n569), .Q(n106) );
  AO22X1 U196 ( .IN1(ctrlFU0_o[9]), .IN2(n571), .IN3(exePacket0_i[82]), .IN4(
        n569), .Q(n107) );
  AO22X1 U197 ( .IN1(ctrlFU0_o[10]), .IN2(n571), .IN3(exePacket0_i[83]), .IN4(
        n570), .Q(n108) );
  AO22X1 U198 ( .IN1(ctrlFU0_o[11]), .IN2(n571), .IN3(exePacket0_i[84]), .IN4(
        n570), .Q(n109) );
  AO22X1 U199 ( .IN1(ctrlFU0_o[12]), .IN2(n571), .IN3(exePacket0_i[85]), .IN4(
        n570), .Q(n110) );
  AO22X1 U200 ( .IN1(ctrlFU0_o[13]), .IN2(n571), .IN3(exePacket0_i[86]), .IN4(
        n570), .Q(n111) );
  AO22X1 U201 ( .IN1(ctrlFU0_o[14]), .IN2(n573), .IN3(exePacket0_i[87]), .IN4(
        n570), .Q(n112) );
  AO22X1 U202 ( .IN1(bypassPacket0_o[35]), .IN2(n573), .IN3(exePacket0_i[88]), 
        .IN4(n570), .Q(n113) );
  AO22X1 U203 ( .IN1(bypassPacket0_o[36]), .IN2(n573), .IN3(exePacket0_i[89]), 
        .IN4(n570), .Q(n114) );
  AO22X1 U204 ( .IN1(bypassPacket0_o[37]), .IN2(n573), .IN3(exePacket0_i[90]), 
        .IN4(n570), .Q(n115) );
  AO22X1 U205 ( .IN1(bypassPacket0_o[38]), .IN2(n573), .IN3(exePacket0_i[91]), 
        .IN4(n570), .Q(n116) );
  AO22X1 U206 ( .IN1(bypassPacket0_o[39]), .IN2(n573), .IN3(exePacket0_i[92]), 
        .IN4(n570), .Q(n117) );
  AO22X1 U207 ( .IN1(bypassPacket0_o[40]), .IN2(n573), .IN3(exePacket0_i[93]), 
        .IN4(n570), .Q(n118) );
  AO22X1 U208 ( .IN1(bypassPacket0_o[41]), .IN2(n573), .IN3(exePacket0_i[94]), 
        .IN4(n570), .Q(n119) );
  AO22X1 U209 ( .IN1(ctrlFU0_o[0]), .IN2(n573), .IN3(exePacket0_i[95]), .IN4(
        n14), .Q(n120) );
  AO22X1 U210 ( .IN1(ctrlFU0_o[1]), .IN2(n573), .IN3(exePacket0_i[96]), .IN4(
        n14), .Q(n121) );
  AO22X1 U211 ( .IN1(ctrlFU0_o[2]), .IN2(n573), .IN3(exePacket0_i[97]), .IN4(
        n14), .Q(n122) );
  AO22X1 U212 ( .IN1(ctrlFU0_o[3]), .IN2(n573), .IN3(exePacket0_i[98]), .IN4(
        n14), .Q(n123) );
  AO22X1 U213 ( .IN1(ctrlFU0_o[4]), .IN2(n573), .IN3(exePacket0_i[99]), .IN4(
        n14), .Q(n124) );
  AO22X1 U214 ( .IN1(ctrlFU0_o[5]), .IN2(n573), .IN3(exePacket0_i[100]), .IN4(
        n14), .Q(n125) );
  AO22X1 U215 ( .IN1(ctrlFU0_o[6]), .IN2(n573), .IN3(exePacket0_i[101]), .IN4(
        n14), .Q(n126) );
  AO22X1 U216 ( .IN1(ctrlFU0_o[7]), .IN2(n573), .IN3(exePacket0_i[102]), .IN4(
        n14), .Q(n127) );
  AO22X1 U217 ( .IN1(ldViolationPacket_i[0]), .IN2(n5), .IN3(
        ldViolationPacket_o[0]), .IN4(n15), .Q(n128) );
  AO22X1 U218 ( .IN1(ldViolationPacket_i[1]), .IN2(n5), .IN3(
        ldViolationPacket_o[1]), .IN4(n15), .Q(n129) );
  AO22X1 U219 ( .IN1(ldViolationPacket_i[2]), .IN2(n5), .IN3(
        ldViolationPacket_o[2]), .IN4(n15), .Q(n130) );
  AO22X1 U220 ( .IN1(ldViolationPacket_i[3]), .IN2(n5), .IN3(
        ldViolationPacket_o[3]), .IN4(n15), .Q(n131) );
  AO22X1 U221 ( .IN1(ldViolationPacket_i[4]), .IN2(n5), .IN3(
        ldViolationPacket_o[4]), .IN4(n15), .Q(n132) );
  AO22X1 U222 ( .IN1(ldViolationPacket_i[5]), .IN2(n5), .IN3(
        ldViolationPacket_o[5]), .IN4(n15), .Q(n133) );
  AO22X1 U223 ( .IN1(ldViolationPacket_i[6]), .IN2(n5), .IN3(
        ldViolationPacket_o[6]), .IN4(n15), .Q(n134) );
  AO22X1 U224 ( .IN1(ldViolationPacket_i[7]), .IN2(n5), .IN3(
        ldViolationPacket_o[7]), .IN4(n15), .Q(n135) );
  AO22X1 U225 ( .IN1(ctrlBrDirection_o), .IN2(n591), .IN3(exePacket2_i_0), 
        .IN4(n587), .Q(n136) );
  AO22X1 U226 ( .IN1(computedAddr2_o[0]), .IN2(n592), .IN3(exePacket2_i_1), 
        .IN4(n586), .Q(n137) );
  AO22X1 U227 ( .IN1(computedAddr2_o[1]), .IN2(n589), .IN3(exePacket2_i_2), 
        .IN4(n585), .Q(n138) );
  AO22X1 U228 ( .IN1(computedAddr2_o[2]), .IN2(n588), .IN3(exePacket2_i_3), 
        .IN4(n584), .Q(n139) );
  AO22X1 U229 ( .IN1(computedAddr2_o[3]), .IN2(n593), .IN3(exePacket2_i_4), 
        .IN4(n8), .Q(n140) );
  AO22X1 U230 ( .IN1(computedAddr2_o[4]), .IN2(n590), .IN3(exePacket2_i_5), 
        .IN4(n587), .Q(n141) );
  AO22X1 U231 ( .IN1(computedAddr2_o[5]), .IN2(n591), .IN3(exePacket2_i_6), 
        .IN4(n586), .Q(n142) );
  AO22X1 U232 ( .IN1(computedAddr2_o[6]), .IN2(n592), .IN3(exePacket2_i_7), 
        .IN4(n585), .Q(n143) );
  AO22X1 U233 ( .IN1(computedAddr2_o[7]), .IN2(n592), .IN3(exePacket2_i_8), 
        .IN4(n584), .Q(n144) );
  AO22X1 U234 ( .IN1(computedAddr2_o[8]), .IN2(n592), .IN3(exePacket2_i_9), 
        .IN4(n587), .Q(n145) );
  AO22X1 U235 ( .IN1(computedAddr2_o[9]), .IN2(n592), .IN3(exePacket2_i_10), 
        .IN4(n586), .Q(n146) );
  AO22X1 U236 ( .IN1(computedAddr2_o[10]), .IN2(n592), .IN3(exePacket2_i_11), 
        .IN4(n585), .Q(n147) );
  AO22X1 U237 ( .IN1(computedAddr2_o[11]), .IN2(n592), .IN3(exePacket2_i_12), 
        .IN4(n584), .Q(n148) );
  AO22X1 U238 ( .IN1(computedAddr2_o[12]), .IN2(n592), .IN3(exePacket2_i_13), 
        .IN4(n8), .Q(n149) );
  AO22X1 U239 ( .IN1(computedAddr2_o[13]), .IN2(n592), .IN3(exePacket2_i_14), 
        .IN4(n8), .Q(n150) );
  AO22X1 U240 ( .IN1(computedAddr2_o[14]), .IN2(n592), .IN3(exePacket2_i_15), 
        .IN4(n8), .Q(n151) );
  AO22X1 U241 ( .IN1(computedAddr2_o[15]), .IN2(n592), .IN3(exePacket2_i_16), 
        .IN4(n8), .Q(n152) );
  AO22X1 U242 ( .IN1(computedAddr2_o[16]), .IN2(n592), .IN3(exePacket2_i_17), 
        .IN4(n587), .Q(n153) );
  AO22X1 U243 ( .IN1(computedAddr2_o[17]), .IN2(n591), .IN3(exePacket2_i_18), 
        .IN4(n587), .Q(n154) );
  AO22X1 U244 ( .IN1(computedAddr2_o[18]), .IN2(n591), .IN3(exePacket2_i_19), 
        .IN4(n587), .Q(n155) );
  AO22X1 U245 ( .IN1(computedAddr2_o[19]), .IN2(n591), .IN3(exePacket2_i_20), 
        .IN4(n587), .Q(n156) );
  AO22X1 U246 ( .IN1(computedAddr2_o[20]), .IN2(n591), .IN3(exePacket2_i_21), 
        .IN4(n587), .Q(n157) );
  AO22X1 U247 ( .IN1(computedAddr2_o[21]), .IN2(n591), .IN3(exePacket2_i_22), 
        .IN4(n587), .Q(n158) );
  AO22X1 U248 ( .IN1(computedAddr2_o[22]), .IN2(n591), .IN3(exePacket2_i_23), 
        .IN4(n587), .Q(n159) );
  AO22X1 U249 ( .IN1(computedAddr2_o[23]), .IN2(n591), .IN3(exePacket2_i_24), 
        .IN4(n587), .Q(n160) );
  AO22X1 U250 ( .IN1(computedAddr2_o[24]), .IN2(n591), .IN3(exePacket2_i_25), 
        .IN4(n587), .Q(n161) );
  AO22X1 U251 ( .IN1(computedAddr2_o[25]), .IN2(n591), .IN3(exePacket2_i_26), 
        .IN4(n587), .Q(n162) );
  AO22X1 U252 ( .IN1(computedAddr2_o[26]), .IN2(n591), .IN3(exePacket2_i_27), 
        .IN4(n587), .Q(n163) );
  AO22X1 U253 ( .IN1(computedAddr2_o[27]), .IN2(n590), .IN3(exePacket2_i_28), 
        .IN4(n587), .Q(n164) );
  AO22X1 U254 ( .IN1(computedAddr2_o[28]), .IN2(n590), .IN3(exePacket2_i_29), 
        .IN4(n586), .Q(n165) );
  AO22X1 U255 ( .IN1(computedAddr2_o[29]), .IN2(n590), .IN3(exePacket2_i_30), 
        .IN4(n586), .Q(n166) );
  AO22X1 U256 ( .IN1(computedAddr2_o[30]), .IN2(n590), .IN3(exePacket2_i_31), 
        .IN4(n586), .Q(n167) );
  AO22X1 U257 ( .IN1(computedAddr2_o[31]), .IN2(n590), .IN3(exePacket2_i_32), 
        .IN4(n586), .Q(n168) );
  AO22X1 U258 ( .IN1(ctrlCtiQueueIndex_o[0]), .IN2(n590), .IN3(exePacket2_i_33), .IN4(n586), .Q(n169) );
  AO22X1 U259 ( .IN1(ctrlCtiQueueIndex_o[1]), .IN2(n590), .IN3(exePacket2_i_34), .IN4(n586), .Q(n170) );
  AO22X1 U260 ( .IN1(ctrlCtiQueueIndex_o[2]), .IN2(n590), .IN3(exePacket2_i_35), .IN4(n586), .Q(n171) );
  AO22X1 U261 ( .IN1(ctrlCtiQueueIndex_o[3]), .IN2(n590), .IN3(exePacket2_i_36), .IN4(n586), .Q(n172) );
  AO22X1 U262 ( .IN1(bypassPacket2_o[1]), .IN2(n590), .IN3(exePacket2_i_37), 
        .IN4(n586), .Q(n173) );
  AO22X1 U263 ( .IN1(bypassPacket2_o[2]), .IN2(n589), .IN3(exePacket2_i_38), 
        .IN4(n586), .Q(n174) );
  AO22X1 U264 ( .IN1(bypassPacket2_o[3]), .IN2(n589), .IN3(exePacket2_i[49]), 
        .IN4(n586), .Q(n175) );
  AO22X1 U265 ( .IN1(bypassPacket2_o[4]), .IN2(n589), .IN3(exePacket2_i[50]), 
        .IN4(n586), .Q(n176) );
  AO22X1 U266 ( .IN1(bypassPacket2_o[5]), .IN2(n589), .IN3(exePacket2_i[51]), 
        .IN4(n585), .Q(n177) );
  AO22X1 U267 ( .IN1(bypassPacket2_o[6]), .IN2(n589), .IN3(exePacket2_i[52]), 
        .IN4(n585), .Q(n178) );
  AO22X1 U268 ( .IN1(bypassPacket2_o[7]), .IN2(n589), .IN3(exePacket2_i[53]), 
        .IN4(n585), .Q(n179) );
  AO22X1 U269 ( .IN1(bypassPacket2_o[8]), .IN2(n589), .IN3(exePacket2_i[54]), 
        .IN4(n585), .Q(n180) );
  AO22X1 U270 ( .IN1(bypassPacket2_o[9]), .IN2(n589), .IN3(exePacket2_i[55]), 
        .IN4(n585), .Q(n181) );
  AO22X1 U271 ( .IN1(bypassPacket2_o[10]), .IN2(n589), .IN3(exePacket2_i[56]), 
        .IN4(n585), .Q(n182) );
  AO22X1 U272 ( .IN1(bypassPacket2_o[11]), .IN2(n589), .IN3(exePacket2_i[57]), 
        .IN4(n585), .Q(n183) );
  AO22X1 U273 ( .IN1(bypassPacket2_o[12]), .IN2(n588), .IN3(exePacket2_i[58]), 
        .IN4(n585), .Q(n184) );
  AO22X1 U274 ( .IN1(bypassPacket2_o[13]), .IN2(n588), .IN3(exePacket2_i[59]), 
        .IN4(n585), .Q(n185) );
  AO22X1 U275 ( .IN1(bypassPacket2_o[14]), .IN2(n588), .IN3(exePacket2_i[60]), 
        .IN4(n585), .Q(n186) );
  AO22X1 U276 ( .IN1(bypassPacket2_o[15]), .IN2(n588), .IN3(exePacket2_i[61]), 
        .IN4(n585), .Q(n187) );
  AO22X1 U277 ( .IN1(bypassPacket2_o[16]), .IN2(n588), .IN3(exePacket2_i[62]), 
        .IN4(n585), .Q(n188) );
  AO22X1 U278 ( .IN1(bypassPacket2_o[17]), .IN2(n588), .IN3(exePacket2_i[63]), 
        .IN4(n584), .Q(n189) );
  AO22X1 U279 ( .IN1(bypassPacket2_o[18]), .IN2(n588), .IN3(exePacket2_i[64]), 
        .IN4(n584), .Q(n190) );
  AO22X1 U280 ( .IN1(bypassPacket2_o[19]), .IN2(n588), .IN3(exePacket2_i[65]), 
        .IN4(n584), .Q(n191) );
  AO22X1 U281 ( .IN1(bypassPacket2_o[20]), .IN2(n588), .IN3(exePacket2_i[66]), 
        .IN4(n584), .Q(n192) );
  AO22X1 U282 ( .IN1(bypassPacket2_o[21]), .IN2(n588), .IN3(exePacket2_i[67]), 
        .IN4(n584), .Q(n193) );
  AO22X1 U283 ( .IN1(bypassPacket2_o[22]), .IN2(n593), .IN3(exePacket2_i[68]), 
        .IN4(n584), .Q(n194) );
  AO22X1 U284 ( .IN1(bypassPacket2_o[23]), .IN2(n590), .IN3(exePacket2_i[69]), 
        .IN4(n584), .Q(n195) );
  AO22X1 U285 ( .IN1(bypassPacket2_o[24]), .IN2(n591), .IN3(exePacket2_i[70]), 
        .IN4(n584), .Q(n196) );
  AO22X1 U286 ( .IN1(bypassPacket2_o[25]), .IN2(n592), .IN3(exePacket2_i[71]), 
        .IN4(n584), .Q(n197) );
  AO22X1 U287 ( .IN1(bypassPacket2_o[26]), .IN2(n589), .IN3(exePacket2_i[72]), 
        .IN4(n584), .Q(n198) );
  AO22X1 U288 ( .IN1(bypassPacket2_o[27]), .IN2(n588), .IN3(exePacket2_i[73]), 
        .IN4(n584), .Q(n199) );
  AO22X1 U289 ( .IN1(bypassPacket2_o[28]), .IN2(n593), .IN3(exePacket2_i[74]), 
        .IN4(n584), .Q(n200) );
  AND2X1 U290 ( .IN1(agenIqFreedValid0_o), .IN2(ctrlFU3_o[4]), .Q(
        bypassValid3_o) );
  AND2X1 U291 ( .IN1(ctrlVerified_o), .IN2(ctrlFU2_o[4]), .Q(bypassValid2_o)
         );
  AND2X1 U292 ( .IN1(exePacketValid1), .IN2(ctrlFU1_o[4]), .Q(bypassValid1_o)
         );
  AND2X1 U293 ( .IN1(exePacketValid0), .IN2(ctrlFU0_o[4]), .Q(bypassValid0_o)
         );
  INVX0 U294 ( .INP(1'b1), .ZN(ctrlMispredict_o) );
  INVX0 U296 ( .INP(1'b1), .ZN(computedAddr3_o[0]) );
  INVX0 U298 ( .INP(1'b1), .ZN(computedAddr3_o[1]) );
  INVX0 U300 ( .INP(1'b1), .ZN(computedAddr3_o[2]) );
  INVX0 U302 ( .INP(1'b1), .ZN(computedAddr3_o[3]) );
  INVX0 U304 ( .INP(1'b1), .ZN(computedAddr3_o[4]) );
  INVX0 U306 ( .INP(1'b1), .ZN(computedAddr3_o[5]) );
  INVX0 U308 ( .INP(1'b1), .ZN(computedAddr3_o[6]) );
  INVX0 U310 ( .INP(1'b1), .ZN(computedAddr3_o[7]) );
  INVX0 U312 ( .INP(1'b1), .ZN(computedAddr3_o[8]) );
  INVX0 U314 ( .INP(1'b1), .ZN(computedAddr3_o[9]) );
  INVX0 U316 ( .INP(1'b1), .ZN(computedAddr3_o[10]) );
  INVX0 U318 ( .INP(1'b1), .ZN(computedAddr3_o[11]) );
  INVX0 U320 ( .INP(1'b1), .ZN(computedAddr3_o[12]) );
  INVX0 U322 ( .INP(1'b1), .ZN(computedAddr3_o[13]) );
  INVX0 U324 ( .INP(1'b1), .ZN(computedAddr3_o[14]) );
  INVX0 U326 ( .INP(1'b1), .ZN(computedAddr3_o[15]) );
  INVX0 U328 ( .INP(1'b1), .ZN(computedAddr3_o[16]) );
  INVX0 U330 ( .INP(1'b1), .ZN(computedAddr3_o[17]) );
  INVX0 U332 ( .INP(1'b1), .ZN(computedAddr3_o[18]) );
  INVX0 U334 ( .INP(1'b1), .ZN(computedAddr3_o[19]) );
  INVX0 U336 ( .INP(1'b1), .ZN(computedAddr3_o[20]) );
  INVX0 U338 ( .INP(1'b1), .ZN(computedAddr3_o[21]) );
  INVX0 U340 ( .INP(1'b1), .ZN(computedAddr3_o[22]) );
  INVX0 U342 ( .INP(1'b1), .ZN(computedAddr3_o[23]) );
  INVX0 U344 ( .INP(1'b1), .ZN(computedAddr3_o[24]) );
  INVX0 U346 ( .INP(1'b1), .ZN(computedAddr3_o[25]) );
  INVX0 U348 ( .INP(1'b1), .ZN(computedAddr3_o[26]) );
  INVX0 U350 ( .INP(1'b1), .ZN(computedAddr3_o[27]) );
  INVX0 U352 ( .INP(1'b1), .ZN(computedAddr3_o[28]) );
  INVX0 U354 ( .INP(1'b1), .ZN(computedAddr3_o[29]) );
  INVX0 U356 ( .INP(1'b1), .ZN(computedAddr3_o[30]) );
  INVX0 U358 ( .INP(1'b1), .ZN(computedAddr3_o[31]) );
  INVX0 U360 ( .INP(1'b1), .ZN(bypassPacket3_o[0]) );
  INVX0 U362 ( .INP(1'b1), .ZN(bypassPacket3_o[1]) );
  INVX0 U364 ( .INP(1'b1), .ZN(bypassPacket3_o[2]) );
  INVX0 U366 ( .INP(1'b1), .ZN(bypassPacket2_o[0]) );
  INVX0 U368 ( .INP(1'b1), .ZN(computedAddr1_o[0]) );
  INVX0 U370 ( .INP(1'b1), .ZN(computedAddr1_o[1]) );
  INVX0 U372 ( .INP(1'b1), .ZN(computedAddr1_o[2]) );
  INVX0 U374 ( .INP(1'b1), .ZN(computedAddr1_o[3]) );
  INVX0 U376 ( .INP(1'b1), .ZN(computedAddr1_o[4]) );
  INVX0 U378 ( .INP(1'b1), .ZN(computedAddr1_o[5]) );
  INVX0 U380 ( .INP(1'b1), .ZN(computedAddr1_o[6]) );
  INVX0 U382 ( .INP(1'b1), .ZN(computedAddr1_o[7]) );
  INVX0 U384 ( .INP(1'b1), .ZN(computedAddr1_o[8]) );
  INVX0 U386 ( .INP(1'b1), .ZN(computedAddr1_o[9]) );
  INVX0 U388 ( .INP(1'b1), .ZN(computedAddr1_o[10]) );
  INVX0 U390 ( .INP(1'b1), .ZN(computedAddr1_o[11]) );
  INVX0 U392 ( .INP(1'b1), .ZN(computedAddr1_o[12]) );
  INVX0 U394 ( .INP(1'b1), .ZN(computedAddr1_o[13]) );
  INVX0 U396 ( .INP(1'b1), .ZN(computedAddr1_o[14]) );
  INVX0 U398 ( .INP(1'b1), .ZN(computedAddr1_o[15]) );
  INVX0 U400 ( .INP(1'b1), .ZN(computedAddr1_o[16]) );
  INVX0 U402 ( .INP(1'b1), .ZN(computedAddr1_o[17]) );
  INVX0 U404 ( .INP(1'b1), .ZN(computedAddr1_o[18]) );
  INVX0 U406 ( .INP(1'b1), .ZN(computedAddr1_o[19]) );
  INVX0 U408 ( .INP(1'b1), .ZN(computedAddr1_o[20]) );
  INVX0 U410 ( .INP(1'b1), .ZN(computedAddr1_o[21]) );
  INVX0 U412 ( .INP(1'b1), .ZN(computedAddr1_o[22]) );
  INVX0 U414 ( .INP(1'b1), .ZN(computedAddr1_o[23]) );
  INVX0 U416 ( .INP(1'b1), .ZN(computedAddr1_o[24]) );
  INVX0 U418 ( .INP(1'b1), .ZN(computedAddr1_o[25]) );
  INVX0 U420 ( .INP(1'b1), .ZN(computedAddr1_o[26]) );
  INVX0 U422 ( .INP(1'b1), .ZN(computedAddr1_o[27]) );
  INVX0 U424 ( .INP(1'b1), .ZN(computedAddr1_o[28]) );
  INVX0 U426 ( .INP(1'b1), .ZN(computedAddr1_o[29]) );
  INVX0 U428 ( .INP(1'b1), .ZN(computedAddr1_o[30]) );
  INVX0 U430 ( .INP(1'b1), .ZN(computedAddr1_o[31]) );
  INVX0 U432 ( .INP(1'b1), .ZN(bypassPacket1_o[0]) );
  INVX0 U434 ( .INP(1'b1), .ZN(computedAddr0_o[0]) );
  INVX0 U436 ( .INP(1'b1), .ZN(computedAddr0_o[1]) );
  INVX0 U438 ( .INP(1'b1), .ZN(computedAddr0_o[2]) );
  INVX0 U440 ( .INP(1'b1), .ZN(computedAddr0_o[3]) );
  INVX0 U442 ( .INP(1'b1), .ZN(computedAddr0_o[4]) );
  INVX0 U444 ( .INP(1'b1), .ZN(computedAddr0_o[5]) );
  INVX0 U446 ( .INP(1'b1), .ZN(computedAddr0_o[6]) );
  INVX0 U448 ( .INP(1'b1), .ZN(computedAddr0_o[7]) );
  INVX0 U450 ( .INP(1'b1), .ZN(computedAddr0_o[8]) );
  INVX0 U452 ( .INP(1'b1), .ZN(computedAddr0_o[9]) );
  INVX0 U454 ( .INP(1'b1), .ZN(computedAddr0_o[10]) );
  INVX0 U456 ( .INP(1'b1), .ZN(computedAddr0_o[11]) );
  INVX0 U458 ( .INP(1'b1), .ZN(computedAddr0_o[12]) );
  INVX0 U460 ( .INP(1'b1), .ZN(computedAddr0_o[13]) );
  INVX0 U462 ( .INP(1'b1), .ZN(computedAddr0_o[14]) );
  INVX0 U464 ( .INP(1'b1), .ZN(computedAddr0_o[15]) );
  INVX0 U466 ( .INP(1'b1), .ZN(computedAddr0_o[16]) );
  INVX0 U468 ( .INP(1'b1), .ZN(computedAddr0_o[17]) );
  INVX0 U470 ( .INP(1'b1), .ZN(computedAddr0_o[18]) );
  INVX0 U472 ( .INP(1'b1), .ZN(computedAddr0_o[19]) );
  INVX0 U474 ( .INP(1'b1), .ZN(computedAddr0_o[20]) );
  INVX0 U476 ( .INP(1'b1), .ZN(computedAddr0_o[21]) );
  INVX0 U478 ( .INP(1'b1), .ZN(computedAddr0_o[22]) );
  INVX0 U480 ( .INP(1'b1), .ZN(computedAddr0_o[23]) );
  INVX0 U482 ( .INP(1'b1), .ZN(computedAddr0_o[24]) );
  INVX0 U484 ( .INP(1'b1), .ZN(computedAddr0_o[25]) );
  INVX0 U486 ( .INP(1'b1), .ZN(computedAddr0_o[26]) );
  INVX0 U488 ( .INP(1'b1), .ZN(computedAddr0_o[27]) );
  INVX0 U490 ( .INP(1'b1), .ZN(computedAddr0_o[28]) );
  INVX0 U492 ( .INP(1'b1), .ZN(computedAddr0_o[29]) );
  INVX0 U494 ( .INP(1'b1), .ZN(computedAddr0_o[30]) );
  INVX0 U496 ( .INP(1'b1), .ZN(computedAddr0_o[31]) );
  INVX0 U498 ( .INP(1'b1), .ZN(bypassPacket0_o[0]) );
  NBUFFX2 U500 ( .INP(n8), .Z(n587) );
  NBUFFX2 U501 ( .INP(n8), .Z(n586) );
  NBUFFX2 U502 ( .INP(n8), .Z(n585) );
  NBUFFX2 U503 ( .INP(n8), .Z(n584) );
  NBUFFX2 U504 ( .INP(n7), .Z(n593) );
  NBUFFX2 U505 ( .INP(n12), .Z(n576) );
  NBUFFX2 U506 ( .INP(n9), .Z(n583) );
  NBUFFX2 U507 ( .INP(n11), .Z(n578) );
  NBUFFX2 U508 ( .INP(n13), .Z(n573) );
  NBUFFX2 U509 ( .INP(n7), .Z(n589) );
  NBUFFX2 U510 ( .INP(n7), .Z(n588) );
  INVX0 U511 ( .INP(n15), .ZN(n5) );
  INVX0 U512 ( .INP(n494), .ZN(ctrlTargetAddr_o[0]) );
  INVX0 U513 ( .INP(n495), .ZN(ctrlTargetAddr_o[1]) );
  INVX0 U514 ( .INP(n496), .ZN(ctrlTargetAddr_o[2]) );
  INVX0 U515 ( .INP(n497), .ZN(ctrlTargetAddr_o[3]) );
  INVX0 U516 ( .INP(n498), .ZN(ctrlTargetAddr_o[4]) );
  INVX0 U517 ( .INP(n499), .ZN(ctrlTargetAddr_o[5]) );
  INVX0 U518 ( .INP(n500), .ZN(ctrlTargetAddr_o[6]) );
  INVX0 U519 ( .INP(n501), .ZN(ctrlTargetAddr_o[7]) );
  INVX0 U520 ( .INP(n502), .ZN(ctrlTargetAddr_o[8]) );
  INVX0 U521 ( .INP(n503), .ZN(ctrlTargetAddr_o[9]) );
  INVX0 U522 ( .INP(n504), .ZN(ctrlTargetAddr_o[10]) );
  INVX0 U523 ( .INP(n505), .ZN(ctrlTargetAddr_o[11]) );
  INVX0 U524 ( .INP(n506), .ZN(ctrlTargetAddr_o[12]) );
  INVX0 U525 ( .INP(n507), .ZN(ctrlTargetAddr_o[13]) );
  NOR2X0 U526 ( .IN1(reset), .IN2(exePacketValid2_i), .QN(n7) );
  NOR2X0 U527 ( .IN1(n7), .IN2(reset), .QN(n8) );
  NOR2X0 U528 ( .IN1(n582), .IN2(reset), .QN(n10) );
  NOR2X0 U529 ( .IN1(n577), .IN2(reset), .QN(n12) );
  NOR2X0 U530 ( .IN1(n13), .IN2(reset), .QN(n14) );
  NOR2X0 U531 ( .IN1(reset), .IN2(exePacketValid1_i), .QN(n11) );
  NOR2X0 U532 ( .IN1(reset), .IN2(exePacketValid0_i), .QN(n13) );
  NOR2X0 U533 ( .IN1(reset), .IN2(lsuPacketValid0_i), .QN(n9) );
  NAND2X1 U534 ( .IN1(lsuPacketValid0_i), .IN2(n6), .QN(n15) );
  INVX0 U535 ( .INP(reset), .ZN(n6) );
  INVX0 U536 ( .INP(n528), .ZN(ctrlConditional_o) );
  INVX0 U537 ( .INP(n527), .ZN(ctrlSMTid_o[1]) );
  INVX0 U538 ( .INP(n526), .ZN(ctrlSMTid_o[0]) );
  INVX0 U539 ( .INP(n563), .ZN(writebkValid3_o) );
  INVX0 U540 ( .INP(n561), .ZN(writebkValid2_o) );
  INVX0 U541 ( .INP(n525), .ZN(ctrlTargetAddr_o[31]) );
  INVX0 U542 ( .INP(n524), .ZN(ctrlTargetAddr_o[30]) );
  INVX0 U543 ( .INP(n523), .ZN(ctrlTargetAddr_o[29]) );
  INVX0 U544 ( .INP(n522), .ZN(ctrlTargetAddr_o[28]) );
  INVX0 U545 ( .INP(n521), .ZN(ctrlTargetAddr_o[27]) );
  INVX0 U546 ( .INP(n520), .ZN(ctrlTargetAddr_o[26]) );
  INVX0 U547 ( .INP(n519), .ZN(ctrlTargetAddr_o[25]) );
  INVX0 U548 ( .INP(n518), .ZN(ctrlTargetAddr_o[24]) );
  INVX0 U549 ( .INP(n517), .ZN(ctrlTargetAddr_o[23]) );
  INVX0 U550 ( .INP(n516), .ZN(ctrlTargetAddr_o[22]) );
  INVX0 U551 ( .INP(n515), .ZN(ctrlTargetAddr_o[21]) );
  INVX0 U552 ( .INP(n514), .ZN(ctrlTargetAddr_o[20]) );
  INVX0 U553 ( .INP(n513), .ZN(ctrlTargetAddr_o[19]) );
  INVX0 U554 ( .INP(n512), .ZN(ctrlTargetAddr_o[18]) );
  INVX0 U555 ( .INP(n511), .ZN(ctrlTargetAddr_o[17]) );
  INVX0 U556 ( .INP(n510), .ZN(ctrlTargetAddr_o[16]) );
  INVX0 U557 ( .INP(n509), .ZN(ctrlTargetAddr_o[15]) );
  INVX0 U558 ( .INP(n508), .ZN(ctrlTargetAddr_o[14]) );
  NBUFFX2 U559 ( .INP(n14), .Z(n568) );
  NBUFFX2 U560 ( .INP(n14), .Z(n569) );
  NBUFFX2 U561 ( .INP(n14), .Z(n570) );
  NBUFFX2 U562 ( .INP(n13), .Z(n571) );
  NBUFFX2 U563 ( .INP(n13), .Z(n572) );
  NBUFFX2 U564 ( .INP(n12), .Z(n574) );
  NBUFFX2 U565 ( .INP(n12), .Z(n575) );
  NBUFFX2 U566 ( .INP(n11), .Z(n577) );
  NBUFFX2 U567 ( .INP(n10), .Z(n579) );
  NBUFFX2 U568 ( .INP(n10), .Z(n580) );
  NBUFFX2 U569 ( .INP(n10), .Z(n581) );
  NBUFFX2 U570 ( .INP(n9), .Z(n582) );
  NBUFFX2 U571 ( .INP(n7), .Z(n590) );
  NBUFFX2 U572 ( .INP(n7), .Z(n591) );
  NBUFFX2 U573 ( .INP(n7), .Z(n592) );
endmodule

