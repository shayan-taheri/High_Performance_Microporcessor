
module Decode_PISA_0 ( instPacketValid_i, instPacket_i, decodedPacket0Valid_o, 
        decodedPacket0_o, decodedPacket1Valid_o, decodedPacket1_o );
  input [132:0] instPacket_i;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  input instPacketValid_i;
  output decodedPacket0Valid_o, decodedPacket1Valid_o;
  wire   instPacket_i_98, instPacket_i_97, instPacket_i_96, instPacket_i_95,
         instPacket_i_94, instPacket_i_93, instPacket_i_92, instPacket_i_91,
         instPacket_i_90, instPacket_i_89, instPacket_i_88, instPacket_i_87,
         instPacket_i_86, instPacket_i_85, instPacket_i_84, instPacket_i_83,
         instPacket_i_82, instPacket_i_81, instPacket_i_80, instPacket_i_79,
         instPacket_i_78, instPacket_i_77, instPacket_i_76, instPacket_i_75,
         instPacket_i_74, instPacket_i_73, instPacket_i_72, instPacket_i_71,
         instPacket_i_36, instPacket_i_35, instPacket_i_34, instPacket_i_33,
         instPacket_i_32, instPacket_i_31, instPacket_i_30, instPacket_i_29,
         instPacket_i_28, instPacket_i_27, instPacket_i_26, instPacket_i_25,
         instPacket_i_24, instPacket_i_23, instPacket_i_22, instPacket_i_21,
         instPacket_i_20, instPacket_i_19, instPacket_i_18, instPacket_i_17,
         instPacket_i_16, instPacket_i_15, instPacket_i_14, instPacket_i_13,
         instPacket_i_12, instPacket_i_11, instPacket_i_10, instPacket_i_9,
         instPacket_i_8, instPacket_i_7, instPacket_i_6, instPacket_i_5, n370,
         decodedPacket1_o_120, decodedPacket1_o_119, decodedPacket1_o_118,
         n371, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         \r340/carry[15] , \r340/carry[14] , \r340/carry[13] ,
         \r340/carry[12] , \r340/carry[11] , \r340/carry[10] , \r340/carry[9] ,
         \r340/carry[8] , \r340/carry[7] , \r340/carry[6] , \r340/carry[5] ,
         \r340/carry[4] , \r339/carry[5] , \r339/carry[4] , \r339/carry[3] ,
         \r339/carry[2] , n306, n307, n311, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369;
  assign instPacket_i_98 = instPacket_i[98];
  assign instPacket_i_97 = instPacket_i[97];
  assign instPacket_i_96 = instPacket_i[96];
  assign instPacket_i_95 = instPacket_i[95];
  assign instPacket_i_94 = instPacket_i[94];
  assign instPacket_i_93 = instPacket_i[93];
  assign instPacket_i_92 = instPacket_i[92];
  assign instPacket_i_91 = instPacket_i[91];
  assign instPacket_i_90 = instPacket_i[90];
  assign instPacket_i_89 = instPacket_i[89];
  assign instPacket_i_88 = instPacket_i[88];
  assign instPacket_i_87 = instPacket_i[87];
  assign instPacket_i_86 = instPacket_i[86];
  assign instPacket_i_85 = instPacket_i[85];
  assign instPacket_i_84 = instPacket_i[84];
  assign instPacket_i_83 = instPacket_i[83];
  assign instPacket_i_82 = instPacket_i[82];
  assign instPacket_i_81 = instPacket_i[81];
  assign instPacket_i_80 = instPacket_i[80];
  assign instPacket_i_79 = instPacket_i[79];
  assign instPacket_i_78 = instPacket_i[78];
  assign instPacket_i_77 = instPacket_i[77];
  assign instPacket_i_76 = instPacket_i[76];
  assign instPacket_i_75 = instPacket_i[75];
  assign instPacket_i_74 = instPacket_i[74];
  assign instPacket_i_73 = instPacket_i[73];
  assign instPacket_i_72 = instPacket_i[72];
  assign instPacket_i_71 = instPacket_i[71];
  assign instPacket_i_36 = instPacket_i[36];
  assign instPacket_i_35 = instPacket_i[35];
  assign instPacket_i_34 = instPacket_i[34];
  assign instPacket_i_33 = instPacket_i[33];
  assign instPacket_i_32 = instPacket_i[32];
  assign instPacket_i_31 = instPacket_i[31];
  assign instPacket_i_30 = instPacket_i[30];
  assign instPacket_i_29 = instPacket_i[29];
  assign instPacket_i_28 = instPacket_i[28];
  assign instPacket_i_27 = instPacket_i[27];
  assign instPacket_i_26 = instPacket_i[26];
  assign instPacket_i_25 = instPacket_i[25];
  assign instPacket_i_24 = instPacket_i[24];
  assign instPacket_i_23 = instPacket_i[23];
  assign instPacket_i_22 = instPacket_i[22];
  assign instPacket_i_21 = instPacket_i[21];
  assign instPacket_i_20 = instPacket_i[20];
  assign instPacket_i_19 = instPacket_i[19];
  assign instPacket_i_18 = instPacket_i[18];
  assign instPacket_i_17 = instPacket_i[17];
  assign instPacket_i_16 = instPacket_i[16];
  assign instPacket_i_15 = instPacket_i[15];
  assign instPacket_i_14 = instPacket_i[14];
  assign instPacket_i_13 = instPacket_i[13];
  assign instPacket_i_12 = instPacket_i[12];
  assign instPacket_i_11 = instPacket_i[11];
  assign instPacket_i_10 = instPacket_i[10];
  assign instPacket_i_9 = instPacket_i[9];
  assign instPacket_i_8 = instPacket_i[8];
  assign instPacket_i_7 = instPacket_i[7];
  assign instPacket_i_6 = instPacket_i[6];
  assign instPacket_i_5 = instPacket_i[5];
  assign decodedPacket1_o[120] = decodedPacket1_o_120;
  assign decodedPacket1_o[119] = decodedPacket1_o_119;
  assign decodedPacket1_o[116] = decodedPacket1_o_118;
  assign N285 = instPacket_i[69];
  assign N286 = instPacket_i[70];

  AND2X1 U160 ( .IN1(N285), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[99]) );
  AO21X1 U161 ( .IN1(N284), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[97]) );
  AND2X1 U162 ( .IN1(decodedPacket1_o_119), .IN2(N283), .Q(
        decodedPacket1_o[96]) );
  AND2X1 U163 ( .IN1(decodedPacket1_o_119), .IN2(N282), .Q(
        decodedPacket1_o[95]) );
  AND2X1 U164 ( .IN1(decodedPacket1_o_119), .IN2(N281), .Q(
        decodedPacket1_o[94]) );
  AND2X1 U165 ( .IN1(decodedPacket1_o_119), .IN2(N280), .Q(
        decodedPacket1_o[93]) );
  AO21X1 U166 ( .IN1(n361), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[92]) );
  OR2X1 U167 ( .IN1(decodedPacket1_o_119), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[91]) );
  AO22X1 U168 ( .IN1(decodedPacket1_o_120), .IN2(N284), .IN3(instPacket_i_90), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[90]) );
  AO22X1 U169 ( .IN1(decodedPacket1_o_120), .IN2(N283), .IN3(instPacket_i_89), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[89]) );
  AO22X1 U170 ( .IN1(decodedPacket1_o_120), .IN2(N282), .IN3(instPacket_i_88), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[88]) );
  AO22X1 U171 ( .IN1(decodedPacket1_o_120), .IN2(N281), .IN3(instPacket_i_87), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[87]) );
  AO22X1 U172 ( .IN1(decodedPacket1_o_120), .IN2(N280), .IN3(instPacket_i_86), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[86]) );
  AO22X1 U173 ( .IN1(decodedPacket1_o_120), .IN2(n361), .IN3(instPacket_i_85), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[85]) );
  OR2X1 U174 ( .IN1(decodedPacket1_o_120), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[84]) );
  AND2X1 U175 ( .IN1(decodedPacket1_o[74]), .IN2(instPacket_i_97), .Q(
        decodedPacket1_o[82]) );
  AND2X1 U176 ( .IN1(decodedPacket1_o[75]), .IN2(instPacket_i_96), .Q(
        decodedPacket1_o[81]) );
  AND2X1 U177 ( .IN1(decodedPacket1_o[73]), .IN2(instPacket_i_95), .Q(
        decodedPacket1_o[80]) );
  AND2X1 U178 ( .IN1(decodedPacket1_o[74]), .IN2(instPacket_i_94), .Q(
        decodedPacket1_o[79]) );
  AND2X1 U179 ( .IN1(N300), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[114]) );
  AND2X1 U180 ( .IN1(N299), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[113]) );
  AND2X1 U181 ( .IN1(N298), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[112]) );
  AND2X1 U182 ( .IN1(N297), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[111]) );
  AND2X1 U183 ( .IN1(N296), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[110]) );
  AND2X1 U184 ( .IN1(N295), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[109]) );
  AND2X1 U185 ( .IN1(N294), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[108]) );
  AND2X1 U186 ( .IN1(N293), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[107]) );
  AND2X1 U187 ( .IN1(N292), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[106]) );
  AND2X1 U188 ( .IN1(N291), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[105]) );
  AND2X1 U189 ( .IN1(N290), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[104]) );
  AND2X1 U190 ( .IN1(N289), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[103]) );
  AND2X1 U191 ( .IN1(N288), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[102]) );
  AND2X1 U192 ( .IN1(N287), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[101]) );
  AND2X1 U193 ( .IN1(N286), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[100]) );
  AND2X1 U194 ( .IN1(instPacketValid_i), .IN2(decodedPacket1_o[73]), .Q(
        decodedPacket1Valid_o) );
  AO22X1 U195 ( .IN1(instPacket_i_9), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_73), .IN4(n311), .Q(decodedPacket0_o[9]) );
  AND2X1 U196 ( .IN1(decodedPacket0_o[98]), .IN2(N285), .Q(
        decodedPacket0_o[99]) );
  AO21X1 U197 ( .IN1(instPacket_i_82), .IN2(n75), .IN3(n76), .Q(n70) );
  OA221X1 U198 ( .IN1(n317), .IN2(n365), .IN3(n74), .IN4(n357), .IN5(n338), 
        .Q(n77) );
  OA221X1 U199 ( .IN1(n317), .IN2(n366), .IN3(n74), .IN4(n358), .IN5(n338), 
        .Q(n78) );
  OA221X1 U200 ( .IN1(n317), .IN2(n367), .IN3(n74), .IN4(n359), .IN5(n338), 
        .Q(n79) );
  OA221X1 U201 ( .IN1(n317), .IN2(n368), .IN3(n74), .IN4(n360), .IN5(n338), 
        .Q(n80) );
  OA221X1 U202 ( .IN1(n317), .IN2(n369), .IN3(n74), .IN4(n361), .IN5(n82), .Q(
        n81) );
  AND3X1 U203 ( .IN1(n84), .IN2(n335), .IN3(n333), .Q(n74) );
  NAND4X0 U204 ( .IN1(n85), .IN2(n318), .IN3(n86), .IN4(n87), .QN(n75) );
  NAND4X0 U205 ( .IN1(n86), .IN2(n338), .IN3(n325), .IN4(n335), .QN(n89) );
  AO22X1 U206 ( .IN1(instPacket_i_8), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_72), .IN4(n67), .Q(decodedPacket0_o[8]) );
  NAND4X0 U207 ( .IN1(n85), .IN2(n330), .IN3(n322), .IN4(n95), .QN(n94) );
  NOR3X0 U208 ( .IN1(n96), .IN2(n332), .IN3(n97), .QN(n95) );
  OA21X1 U209 ( .IN1(n344), .IN2(n345), .IN3(n336), .Q(n96) );
  AND3X1 U210 ( .IN1(n98), .IN2(n319), .IN3(n326), .Q(n85) );
  OA221X1 U211 ( .IN1(n316), .IN2(n354), .IN3(n356), .IN4(n101), .IN5(n102), 
        .Q(n100) );
  AO22X1 U212 ( .IN1(n103), .IN2(instPacket_i_97), .IN3(n104), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[82]) );
  AO22X1 U213 ( .IN1(n103), .IN2(instPacket_i_96), .IN3(n104), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[81]) );
  AO22X1 U214 ( .IN1(n103), .IN2(instPacket_i_95), .IN3(n104), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[80]) );
  AO22X1 U215 ( .IN1(instPacket_i_7), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_71), .IN4(n67), .Q(decodedPacket0_o[7]) );
  AO22X1 U216 ( .IN1(n103), .IN2(instPacket_i_94), .IN3(n104), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[79]) );
  OA221X1 U217 ( .IN1(n316), .IN2(n355), .IN3(n361), .IN4(n101), .IN5(n106), 
        .Q(n105) );
  OA21X1 U218 ( .IN1(n108), .IN2(n107), .IN3(n313), .Q(decodedPacket0_o[77])
         );
  NAND4X0 U219 ( .IN1(n109), .IN2(n326), .IN3(n322), .IN4(n110), .QN(n107) );
  NAND3X0 U220 ( .IN1(n114), .IN2(n87), .IN3(n115), .QN(n90) );
  AO21X1 U221 ( .IN1(instPacket_i[104]), .IN2(n117), .IN3(decodedPacket1_o[72]), .Q(decodedPacket0_o[72]) );
  NAND3X0 U222 ( .IN1(n119), .IN2(n114), .IN3(n120), .QN(n118) );
  AO21X1 U223 ( .IN1(instPacket_i[102]), .IN2(n117), .IN3(decodedPacket1_o[70]), .Q(decodedPacket0_o[70]) );
  AO21X1 U224 ( .IN1(n313), .IN2(n320), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket1_o[70]) );
  AO22X1 U225 ( .IN1(instPacket_i_6), .IN2(decodedPacket0_o[121]), .IN3(N286), 
        .IN4(n67), .Q(decodedPacket0_o[6]) );
  AND2X1 U226 ( .IN1(n117), .IN2(instPacket_i[101]), .Q(decodedPacket0_o[69])
         );
  NAND4X0 U227 ( .IN1(n87), .IN2(n328), .IN3(n121), .IN4(n122), .QN(n117) );
  AND2X1 U228 ( .IN1(instPacket_i[106]), .IN2(n124), .Q(n123) );
  NAND4X0 U229 ( .IN1(n346), .IN2(n339), .IN3(n125), .IN4(n126), .QN(n124) );
  OA22X1 U230 ( .IN1(instPacket_i[105]), .IN2(n351), .IN3(n127), .IN4(n341), 
        .Q(n126) );
  AO22X1 U231 ( .IN1(n99), .IN2(n129), .IN3(n130), .IN4(n131), .Q(n91) );
  NAND4X0 U232 ( .IN1(n133), .IN2(n134), .IN3(n135), .IN4(n136), .QN(n129) );
  NOR3X0 U233 ( .IN1(n137), .IN2(n347), .IN3(n348), .QN(n136) );
  OA21X1 U234 ( .IN1(instPacket_i[103]), .IN2(n125), .IN3(n139), .Q(n138) );
  NAND4X0 U235 ( .IN1(n109), .IN2(n318), .IN3(n140), .IN4(n333), .QN(n92) );
  AND2X1 U236 ( .IN1(n319), .IN2(n141), .Q(n140) );
  OA21X1 U237 ( .IN1(n347), .IN2(n348), .IN3(n324), .Q(n112) );
  AND2X1 U238 ( .IN1(n106), .IN2(n142), .Q(n102) );
  NAND3X0 U239 ( .IN1(n324), .IN2(n353), .IN3(n350), .QN(n142) );
  OR2X1 U240 ( .IN1(n135), .IN2(n132), .Q(n106) );
  AND4X1 U241 ( .IN1(n143), .IN2(n144), .IN3(n145), .IN4(n146), .Q(n109) );
  NOR3X0 U242 ( .IN1(n125), .IN2(instPacket_i[103]), .IN3(n148), .QN(n72) );
  AOI22X1 U243 ( .IN1(n339), .IN2(n340), .IN3(instPacket_i[103]), .IN4(
        instPacket_i[104]), .QN(n121) );
  OR2X1 U244 ( .IN1(n132), .IN2(n149), .Q(n87) );
  AO22X1 U245 ( .IN1(instPacket_i_5), .IN2(decodedPacket0_o[121]), .IN3(N285), 
        .IN4(n67), .Q(decodedPacket0_o[5]) );
  AND2X1 U246 ( .IN1(instPacket_i_36), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[36]) );
  AND2X1 U247 ( .IN1(instPacket_i_35), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[35]) );
  AND2X1 U248 ( .IN1(instPacket_i_34), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[34]) );
  AND2X1 U249 ( .IN1(instPacket_i_33), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[33]) );
  AND2X1 U250 ( .IN1(instPacket_i_32), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[32]) );
  AND2X1 U251 ( .IN1(instPacket_i_31), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[31]) );
  AO22X1 U252 ( .IN1(instPacket_i_30), .IN2(decodedPacket0_o[121]), .IN3(n67), 
        .IN4(instPacket_i_94), .Q(decodedPacket0_o[30]) );
  AO22X1 U253 ( .IN1(instPacket_i_29), .IN2(decodedPacket0_o[121]), .IN3(n67), 
        .IN4(instPacket_i_93), .Q(decodedPacket0_o[29]) );
  AO22X1 U254 ( .IN1(instPacket_i_28), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_92), .IN4(n67), .Q(decodedPacket0_o[28]) );
  AO22X1 U255 ( .IN1(instPacket_i_27), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_91), .IN4(n67), .Q(decodedPacket0_o[27]) );
  AO22X1 U256 ( .IN1(instPacket_i_26), .IN2(n370), .IN3(n67), .IN4(
        instPacket_i_90), .Q(decodedPacket0_o[26]) );
  AO22X1 U257 ( .IN1(instPacket_i_25), .IN2(n370), .IN3(n311), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[25]) );
  AO22X1 U258 ( .IN1(instPacket_i_24), .IN2(n370), .IN3(n67), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[24]) );
  AO22X1 U259 ( .IN1(instPacket_i_23), .IN2(n370), .IN3(n311), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[23]) );
  AO22X1 U260 ( .IN1(instPacket_i_22), .IN2(n370), .IN3(n67), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[22]) );
  AO22X1 U261 ( .IN1(instPacket_i_21), .IN2(n370), .IN3(n67), .IN4(
        instPacket_i_85), .Q(decodedPacket0_o[21]) );
  AO22X1 U262 ( .IN1(instPacket_i_20), .IN2(n370), .IN3(instPacket_i_84), 
        .IN4(n311), .Q(decodedPacket0_o[20]) );
  AO22X1 U263 ( .IN1(instPacket_i_19), .IN2(n370), .IN3(instPacket_i_83), 
        .IN4(n311), .Q(decodedPacket0_o[19]) );
  AO22X1 U264 ( .IN1(instPacket_i_18), .IN2(n370), .IN3(instPacket_i_82), 
        .IN4(n311), .Q(decodedPacket0_o[18]) );
  AO22X1 U265 ( .IN1(instPacket_i_17), .IN2(n370), .IN3(instPacket_i_81), 
        .IN4(n311), .Q(decodedPacket0_o[17]) );
  AO22X1 U266 ( .IN1(instPacket_i_16), .IN2(n370), .IN3(instPacket_i_80), 
        .IN4(n311), .Q(decodedPacket0_o[16]) );
  AO22X1 U267 ( .IN1(instPacket_i_15), .IN2(n370), .IN3(instPacket_i_79), 
        .IN4(n311), .Q(decodedPacket0_o[15]) );
  AO22X1 U268 ( .IN1(instPacket_i_14), .IN2(n370), .IN3(instPacket_i_78), 
        .IN4(n311), .Q(decodedPacket0_o[14]) );
  AO22X1 U269 ( .IN1(instPacket_i_13), .IN2(n370), .IN3(instPacket_i_77), 
        .IN4(n311), .Q(decodedPacket0_o[13]) );
  AO22X1 U270 ( .IN1(instPacket_i_12), .IN2(n370), .IN3(instPacket_i_76), 
        .IN4(n311), .Q(decodedPacket0_o[12]) );
  AO21X1 U271 ( .IN1(n313), .IN2(n150), .IN3(decodedPacket1_o_120), .Q(
        decodedPacket0_o[120]) );
  AO22X1 U272 ( .IN1(instPacket_i_11), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_75), .IN4(n311), .Q(decodedPacket0_o[11]) );
  AO21X1 U273 ( .IN1(n313), .IN2(n152), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket0_o[119]) );
  AO21X1 U274 ( .IN1(n334), .IN2(n155), .IN3(n307), .Q(n154) );
  NOR3X0 U275 ( .IN1(n157), .IN2(n331), .IN3(n158), .QN(n156) );
  NAND3X0 U276 ( .IN1(n163), .IN2(n337), .IN3(n120), .QN(n161) );
  NAND3X0 U277 ( .IN1(n149), .IN2(n166), .IN3(n167), .QN(n165) );
  AND2X1 U278 ( .IN1(n313), .IN2(n168), .Q(decodedPacket0_o[115]) );
  NAND4X0 U279 ( .IN1(n116), .IN2(n333), .IN3(n330), .IN4(n169), .QN(n168) );
  NAND4X0 U280 ( .IN1(n348), .IN2(instPacket_i[106]), .IN3(n341), .IN4(n339), 
        .QN(n169) );
  AND2X1 U281 ( .IN1(n120), .IN2(n321), .Q(n116) );
  NAND3X0 U282 ( .IN1(n325), .IN2(n114), .IN3(n115), .QN(n76) );
  OA21X1 U283 ( .IN1(n134), .IN2(n132), .IN3(n119), .Q(n115) );
  OR2X1 U284 ( .IN1(n132), .IN2(n172), .Q(n114) );
  AO22X1 U285 ( .IN1(instPacket_i_10), .IN2(n370), .IN3(instPacket_i_74), 
        .IN4(n311), .Q(decodedPacket0_o[10]) );
  AND2X1 U286 ( .IN1(n313), .IN2(n162), .Q(n67) );
  AO21X1 U287 ( .IN1(n336), .IN2(n175), .IN3(n83), .Q(n162) );
  OA21X1 U288 ( .IN1(n111), .IN2(n164), .IN3(n313), .Q(n370) );
  AND2X1 U289 ( .IN1(n336), .IN2(n178), .Q(n111) );
  NAND4X0 U290 ( .IN1(n149), .IN2(n147), .IN3(n179), .IN4(n172), .QN(n178) );
  AND2X1 U291 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_76), .Q(
        decodedPacket0_o[106]) );
  AND2X1 U292 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_75), .Q(
        decodedPacket0_o[105]) );
  AND2X1 U293 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_74), .Q(
        decodedPacket0_o[104]) );
  AND2X1 U294 ( .IN1(instPacket_i_73), .IN2(decodedPacket0_o[98]), .Q(
        decodedPacket0_o[103]) );
  AND2X1 U295 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_72), .Q(
        decodedPacket0_o[102]) );
  AND2X1 U296 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_71), .Q(
        decodedPacket0_o[101]) );
  AND2X1 U297 ( .IN1(decodedPacket0_o[98]), .IN2(N286), .Q(
        decodedPacket0_o[100]) );
  OA21X1 U298 ( .IN1(n181), .IN2(n327), .IN3(n313), .Q(decodedPacket0_o[98])
         );
  NAND4X0 U299 ( .IN1(n182), .IN2(n183), .IN3(n184), .IN4(n185), .QN(n69) );
  OR3X1 U300 ( .IN1(instPacket_i[132]), .IN2(instPacket_i[131]), .IN3(
        instPacket_i[130]), .Q(n186) );
  OR3X1 U301 ( .IN1(instPacket_i[126]), .IN2(instPacket_i[125]), .IN3(
        instPacket_i[124]), .Q(n187) );
  OR3X1 U302 ( .IN1(instPacket_i[120]), .IN2(instPacket_i[119]), .IN3(
        instPacket_i[118]), .Q(n188) );
  OR3X1 U303 ( .IN1(instPacket_i[114]), .IN2(instPacket_i[113]), .IN3(
        instPacket_i[112]), .Q(n189) );
  NAND3X0 U304 ( .IN1(n173), .IN2(n191), .IN3(n172), .QN(n190) );
  NAND3X0 U305 ( .IN1(n329), .IN2(n192), .IN3(n84), .QN(n181) );
  AND4X1 U306 ( .IN1(n143), .IN2(n144), .IN3(n193), .IN4(n141), .Q(n84) );
  NAND4X0 U307 ( .IN1(n347), .IN2(instPacket_i[106]), .IN3(n341), .IN4(n339), 
        .QN(n141) );
  AOI22X1 U308 ( .IN1(n175), .IN2(n324), .IN3(n99), .IN4(n194), .QN(n144) );
  AO22X1 U309 ( .IN1(n350), .IN2(n353), .IN3(n131), .IN4(instPacket_i[103]), 
        .Q(n194) );
  NAND3X0 U310 ( .IN1(instPacket_i[103]), .IN2(n352), .IN3(instPacket_i[104]), 
        .QN(n139) );
  AOI222X1 U311 ( .IN1(n99), .IN2(n175), .IN3(n195), .IN4(n323), .IN5(n349), 
        .IN6(n324), .QN(n143) );
  NAND3X0 U312 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[101]), .IN3(n128), 
        .QN(n166) );
  AND3X1 U313 ( .IN1(instPacket_i[101]), .IN2(n352), .IN3(n128), .Q(n175) );
  AND2X1 U314 ( .IN1(n196), .IN2(instPacket_i[105]), .Q(n99) );
  AND3X1 U315 ( .IN1(n340), .IN2(n328), .IN3(instPacket_i[107]), .Q(n196) );
  AO21X1 U316 ( .IN1(n167), .IN2(n191), .IN3(n177), .Q(n192) );
  AND3X1 U317 ( .IN1(n180), .IN2(n172), .IN3(n179), .Q(n167) );
  AND2X1 U318 ( .IN1(n134), .IN2(n173), .Q(n179) );
  NAND3X0 U319 ( .IN1(instPacket_i[101]), .IN2(n197), .IN3(instPacket_i[102]), 
        .QN(n172) );
  NAND4X0 U320 ( .IN1(n330), .IN2(n170), .IN3(n198), .IN4(n120), .QN(n113) );
  NAND3X0 U321 ( .IN1(n197), .IN2(n352), .IN3(instPacket_i[101]), .QN(n191) );
  AND3X1 U322 ( .IN1(n352), .IN2(n351), .IN3(instPacket_i[104]), .Q(n201) );
  NAND3X0 U323 ( .IN1(n341), .IN2(n340), .IN3(n202), .QN(n177) );
  NOR3X0 U324 ( .IN1(n157), .IN2(n158), .IN3(n203), .QN(n170) );
  AOI21X1 U325 ( .IN1(n176), .IN2(n204), .IN3(n200), .QN(n203) );
  NAND3X0 U326 ( .IN1(n202), .IN2(n341), .IN3(instPacket_i[106]), .QN(n200) );
  NAND3X0 U327 ( .IN1(n197), .IN2(n353), .IN3(instPacket_i[102]), .QN(n180) );
  NAND3X0 U328 ( .IN1(n155), .IN2(n159), .IN3(n205), .QN(n150) );
  NAND3X0 U329 ( .IN1(n353), .IN2(n352), .IN3(n128), .QN(n204) );
  NAND3X0 U330 ( .IN1(instPacket_i[102]), .IN2(n353), .IN3(n128), .QN(n176) );
  AND3X1 U331 ( .IN1(instPacket_i[105]), .IN2(n202), .IN3(instPacket_i[106]), 
        .Q(n199) );
  NAND3X0 U332 ( .IN1(n353), .IN2(n352), .IN3(n197), .QN(n133) );
  HADDX1 \r339/U1_1_1  ( .A0(instPacket_i_86), .B0(instPacket_i_85), .C1(
        \r339/carry[2] ), .SO(N280) );
  HADDX1 \r339/U1_1_2  ( .A0(instPacket_i_87), .B0(\r339/carry[2] ), .C1(
        \r339/carry[3] ), .SO(N281) );
  HADDX1 \r339/U1_1_3  ( .A0(instPacket_i_88), .B0(\r339/carry[3] ), .C1(
        \r339/carry[4] ), .SO(N282) );
  HADDX1 \r339/U1_1_4  ( .A0(instPacket_i_89), .B0(\r339/carry[4] ), .C1(
        \r339/carry[5] ), .SO(N283) );
  INVX0 U3 ( .INP(1'b1), .ZN(decodedPacket1_o[5]) );
  INVX0 U5 ( .INP(1'b1), .ZN(decodedPacket1_o[6]) );
  INVX0 U7 ( .INP(1'b1), .ZN(decodedPacket1_o[7]) );
  INVX0 U9 ( .INP(1'b1), .ZN(decodedPacket1_o[8]) );
  INVX0 U11 ( .INP(1'b1), .ZN(decodedPacket1_o[9]) );
  INVX0 U13 ( .INP(1'b1), .ZN(decodedPacket1_o[10]) );
  INVX0 U15 ( .INP(1'b1), .ZN(decodedPacket1_o[11]) );
  INVX0 U17 ( .INP(1'b1), .ZN(decodedPacket1_o[12]) );
  INVX0 U19 ( .INP(1'b1), .ZN(decodedPacket1_o[13]) );
  INVX0 U21 ( .INP(1'b1), .ZN(decodedPacket1_o[14]) );
  INVX0 U23 ( .INP(1'b1), .ZN(decodedPacket1_o[15]) );
  INVX0 U25 ( .INP(1'b1), .ZN(decodedPacket1_o[16]) );
  INVX0 U27 ( .INP(1'b1), .ZN(decodedPacket1_o[17]) );
  INVX0 U29 ( .INP(1'b1), .ZN(decodedPacket1_o[18]) );
  INVX0 U31 ( .INP(1'b1), .ZN(decodedPacket1_o[19]) );
  INVX0 U33 ( .INP(1'b1), .ZN(decodedPacket1_o[20]) );
  INVX0 U35 ( .INP(1'b1), .ZN(decodedPacket1_o[21]) );
  INVX0 U37 ( .INP(1'b1), .ZN(decodedPacket1_o[22]) );
  INVX0 U39 ( .INP(1'b1), .ZN(decodedPacket1_o[23]) );
  INVX0 U41 ( .INP(1'b1), .ZN(decodedPacket1_o[24]) );
  INVX0 U43 ( .INP(1'b1), .ZN(decodedPacket1_o[25]) );
  INVX0 U45 ( .INP(1'b1), .ZN(decodedPacket1_o[26]) );
  INVX0 U47 ( .INP(1'b1), .ZN(decodedPacket1_o[27]) );
  INVX0 U49 ( .INP(1'b1), .ZN(decodedPacket1_o[28]) );
  INVX0 U51 ( .INP(1'b1), .ZN(decodedPacket1_o[29]) );
  INVX0 U53 ( .INP(1'b1), .ZN(decodedPacket1_o[30]) );
  INVX0 U55 ( .INP(1'b1), .ZN(decodedPacket1_o[31]) );
  INVX0 U57 ( .INP(1'b1), .ZN(decodedPacket1_o[32]) );
  INVX0 U59 ( .INP(1'b1), .ZN(decodedPacket1_o[33]) );
  INVX0 U61 ( .INP(1'b1), .ZN(decodedPacket1_o[34]) );
  INVX0 U63 ( .INP(1'b1), .ZN(decodedPacket1_o[35]) );
  INVX0 U65 ( .INP(1'b1), .ZN(decodedPacket1_o[36]) );
  INVX0 U67 ( .INP(1'b1), .ZN(decodedPacket1_o[117]) );
  INVX0 U69 ( .INP(1'b1), .ZN(decodedPacket1_o[121]) );
  INVX0 U71 ( .INP(1'b1), .ZN(decodedPacket1_o[122]) );
  INVX0 U73 ( .INP(1'b1), .ZN(decodedPacket1_o[123]) );
  INVX0 U75 ( .INP(1'b1), .ZN(decodedPacket1_o[124]) );
  INVX0 U77 ( .INP(1'b1), .ZN(decodedPacket1_o[125]) );
  INVX0 U79 ( .INP(1'b1), .ZN(decodedPacket0_o[122]) );
  INVX0 U81 ( .INP(1'b1), .ZN(decodedPacket0_o[123]) );
  INVX0 U83 ( .INP(1'b1), .ZN(decodedPacket0_o[124]) );
  INVX0 U85 ( .INP(1'b1), .ZN(decodedPacket0_o[125]) );
  INVX0 U87 ( .INP(decodedPacket1_o[74]), .ZN(n315) );
  NBUFFX2 U88 ( .INP(decodedPacket1_o[75]), .Z(decodedPacket1_o[69]) );
  NBUFFX2 U89 ( .INP(decodedPacket1_o[75]), .Z(decodedPacket1_o[115]) );
  NBUFFX2 U90 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[77]) );
  NBUFFX2 U91 ( .INP(decodedPacket1_o[73]), .Z(decodedPacket1_o[76]) );
  NBUFFX2 U92 ( .INP(n371), .Z(decodedPacket1_o[73]) );
  NBUFFX2 U93 ( .INP(n371), .Z(decodedPacket1_o[75]) );
  NBUFFX2 U94 ( .INP(n371), .Z(decodedPacket1_o[74]) );
  INVX0 U95 ( .INP(decodedPacket1_o[98]), .ZN(n314) );
  NBUFFX2 U96 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[98]) );
  NBUFFX2 U97 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[118]) );
  NOR2X0 U98 ( .IN1(n69), .IN2(n116), .QN(n371) );
  INVX0 U99 ( .INP(n76), .ZN(n321) );
  NOR2X0 U100 ( .IN1(n335), .IN2(n307), .QN(decodedPacket1_o_119) );
  INVX0 U101 ( .INP(n107), .ZN(n316) );
  INVX0 U102 ( .INP(n75), .ZN(n317) );
  NOR2X0 U103 ( .IN1(n307), .IN2(n316), .QN(n103) );
  INVX0 U104 ( .INP(n93), .ZN(decodedPacket0_o[84]) );
  NOR2X0 U105 ( .IN1(n88), .IN2(n306), .QN(decodedPacket0_o[91]) );
  INVX0 U106 ( .INP(n115), .ZN(n320) );
  NAND2X1 U107 ( .IN1(n342), .IN2(n336), .QN(n86) );
  INVX0 U108 ( .INP(n152), .ZN(n333) );
  INVX0 U109 ( .INP(n90), .ZN(n322) );
  NAND2X1 U110 ( .IN1(n314), .IN2(n154), .QN(decodedPacket0_o[118]) );
  INVX0 U111 ( .INP(n66), .ZN(decodedPacket1_o[71]) );
  INVX0 U112 ( .INP(n108), .ZN(n318) );
  INVX0 U113 ( .INP(n112), .ZN(n319) );
  NOR2X0 U114 ( .IN1(n153), .IN2(n332), .QN(n120) );
  INVX0 U115 ( .INP(n151), .ZN(n332) );
  NAND2X1 U116 ( .IN1(n344), .IN2(n324), .QN(n119) );
  INVX0 U117 ( .INP(n132), .ZN(n324) );
  INVX0 U118 ( .INP(n97), .ZN(n325) );
  NOR2X0 U119 ( .IN1(n306), .IN2(n321), .QN(decodedPacket1_o[72]) );
  NOR2X0 U120 ( .IN1(n307), .IN2(n120), .QN(decodedPacket1_o_118) );
  NAND2X1 U121 ( .IN1(n313), .IN2(n181), .QN(n174) );
  NAND2X1 U122 ( .IN1(n313), .IN2(n94), .QN(n93) );
  INVX0 U123 ( .INP(n69), .ZN(n313) );
  NOR2X0 U124 ( .IN1(n164), .IN2(n171), .QN(n198) );
  NOR2X0 U125 ( .IN1(n156), .IN2(n306), .QN(decodedPacket0_o[117]) );
  INVX0 U126 ( .INP(n159), .ZN(n331) );
  NOR4X0 U127 ( .IN1(n111), .IN2(n112), .IN3(n97), .IN4(n113), .QN(n110) );
  INVX0 U128 ( .INP(n177), .ZN(n336) );
  NOR2X0 U129 ( .IN1(n306), .IN2(n151), .QN(decodedPacket1_o_120) );
  INVX0 U130 ( .INP(n133), .ZN(n342) );
  NOR2X0 U131 ( .IN1(n135), .IN2(n177), .QN(n164) );
  INVX0 U132 ( .INP(n101), .ZN(n327) );
  INVX0 U133 ( .INP(n204), .ZN(n348) );
  INVX0 U134 ( .INP(n153), .ZN(n335) );
  NOR2X0 U135 ( .IN1(n101), .IN2(n307), .QN(n104) );
  NOR2X0 U136 ( .IN1(n342), .IN2(n345), .QN(n149) );
  NAND2X1 U137 ( .IN1(n170), .IN2(n334), .QN(n152) );
  INVX0 U138 ( .INP(n171), .ZN(n334) );
  INVX0 U139 ( .INP(n83), .ZN(n338) );
  NAND2X1 U140 ( .IN1(n313), .IN2(n118), .QN(n66) );
  NOR2X0 U141 ( .IN1(n349), .IN2(n344), .QN(n147) );
  NOR2X0 U142 ( .IN1(n105), .IN2(n307), .QN(decodedPacket0_o[78]) );
  NOR2X0 U143 ( .IN1(n100), .IN2(n306), .QN(decodedPacket0_o[83]) );
  NOR2X0 U144 ( .IN1(n81), .IN2(n307), .QN(decodedPacket0_o[92]) );
  NOR2X0 U145 ( .IN1(n80), .IN2(n307), .QN(decodedPacket0_o[93]) );
  NOR2X0 U146 ( .IN1(n79), .IN2(n307), .QN(decodedPacket0_o[94]) );
  NOR2X0 U147 ( .IN1(n78), .IN2(n306), .QN(decodedPacket0_o[95]) );
  NOR2X0 U148 ( .IN1(n77), .IN2(n306), .QN(decodedPacket0_o[96]) );
  INVX0 U149 ( .INP(n150), .ZN(n330) );
  NAND2X1 U150 ( .IN1(n102), .IN2(n101), .QN(n108) );
  NOR4X0 U151 ( .IN1(n161), .IN2(n162), .IN3(n150), .IN4(n152), .QN(n160) );
  INVX0 U152 ( .INP(n164), .ZN(n337) );
  NAND2X1 U153 ( .IN1(n336), .IN2(n165), .QN(n163) );
  NOR4X0 U154 ( .IN1(n89), .IN2(n90), .IN3(n91), .IN4(n92), .QN(n88) );
  NOR2X0 U155 ( .IN1(n160), .IN2(n307), .QN(decodedPacket0_o[116]) );
  INVX0 U156 ( .INP(n91), .ZN(n326) );
  INVX0 U157 ( .INP(n180), .ZN(n344) );
  INVX0 U158 ( .INP(n191), .ZN(n345) );
  NAND2X1 U159 ( .IN1(n345), .IN2(n199), .QN(n151) );
  NOR2X0 U333 ( .IN1(n173), .IN2(n200), .QN(n153) );
  NAND2X1 U334 ( .IN1(n196), .IN2(n341), .QN(n132) );
  NOR2X0 U335 ( .IN1(n132), .IN2(n173), .QN(n97) );
  NAND2X1 U336 ( .IN1(n201), .IN2(n353), .QN(n134) );
  NAND2X1 U337 ( .IN1(n348), .IN2(n199), .QN(n205) );
  INVX0 U338 ( .INP(n113), .ZN(n329) );
  NOR2X0 U339 ( .IN1(n134), .IN2(n200), .QN(n171) );
  NOR2X0 U340 ( .IN1(n133), .IN2(n200), .QN(n158) );
  NOR2X0 U341 ( .IN1(n180), .IN2(n200), .QN(n157) );
  NOR2X0 U342 ( .IN1(n176), .IN2(n177), .QN(n83) );
  NAND2X1 U343 ( .IN1(n99), .IN2(n190), .QN(n101) );
  INVX0 U344 ( .INP(n176), .ZN(n347) );
  NOR2X0 U345 ( .IN1(n139), .IN2(n148), .QN(n73) );
  INVX0 U346 ( .INP(n166), .ZN(n349) );
  NOR2X0 U347 ( .IN1(n351), .IN2(n132), .QN(n130) );
  NAND2X1 U348 ( .IN1(n131), .IN2(n351), .QN(n135) );
  NAND2X1 U349 ( .IN1(n347), .IN2(n199), .QN(n159) );
  NOR2X0 U350 ( .IN1(n83), .IN2(n72), .QN(n82) );
  NOR2X0 U351 ( .IN1(n315), .IN2(n355), .QN(decodedPacket1_o[78]) );
  NOR2X0 U352 ( .IN1(n315), .IN2(n354), .QN(decodedPacket1_o[83]) );
  NAND2X1 U353 ( .IN1(n66), .IN2(n351), .QN(decodedPacket0_o[71]) );
  NAND2X1 U354 ( .IN1(n315), .IN2(n341), .QN(decodedPacket0_o[73]) );
  NAND2X1 U355 ( .IN1(n315), .IN2(n340), .QN(decodedPacket0_o[74]) );
  NAND2X1 U356 ( .IN1(n315), .IN2(n339), .QN(decodedPacket0_o[75]) );
  NAND2X1 U357 ( .IN1(n315), .IN2(n328), .QN(decodedPacket0_o[76]) );
  NOR2X0 U358 ( .IN1(n361), .IN2(n93), .QN(decodedPacket0_o[85]) );
  NOR2X0 U359 ( .IN1(n360), .IN2(n93), .QN(decodedPacket0_o[86]) );
  NOR2X0 U360 ( .IN1(n359), .IN2(n93), .QN(decodedPacket0_o[87]) );
  NOR2X0 U361 ( .IN1(n358), .IN2(n93), .QN(decodedPacket0_o[88]) );
  NOR2X0 U362 ( .IN1(n357), .IN2(n93), .QN(decodedPacket0_o[89]) );
  NOR2X0 U363 ( .IN1(n356), .IN2(n93), .QN(decodedPacket0_o[90]) );
  NOR2X0 U364 ( .IN1(n68), .IN2(n306), .QN(decodedPacket0_o[97]) );
  NAND2X1 U365 ( .IN1(n342), .IN2(n199), .QN(n155) );
  NAND2X1 U366 ( .IN1(n99), .IN2(n343), .QN(n146) );
  NOR2X0 U367 ( .IN1(n72), .IN2(n73), .QN(n145) );
  INVX0 U368 ( .INP(n147), .ZN(n343) );
  NAND2X1 U369 ( .IN1(n349), .IN2(n99), .QN(n193) );
  NAND2X1 U370 ( .IN1(n99), .IN2(n344), .QN(n98) );
  INVX0 U371 ( .INP(n139), .ZN(n350) );
  NOR2X0 U372 ( .IN1(n369), .IN2(n174), .QN(decodedPacket0_o[107]) );
  NOR2X0 U373 ( .IN1(n368), .IN2(n174), .QN(decodedPacket0_o[108]) );
  NOR2X0 U374 ( .IN1(n367), .IN2(n174), .QN(decodedPacket0_o[109]) );
  NOR2X0 U375 ( .IN1(n366), .IN2(n174), .QN(decodedPacket0_o[110]) );
  NOR2X0 U376 ( .IN1(n365), .IN2(n174), .QN(decodedPacket0_o[111]) );
  NOR2X0 U377 ( .IN1(n364), .IN2(n174), .QN(decodedPacket0_o[112]) );
  NOR2X0 U378 ( .IN1(n363), .IN2(n174), .QN(decodedPacket0_o[113]) );
  NOR2X0 U379 ( .IN1(n362), .IN2(n174), .QN(decodedPacket0_o[114]) );
  INVX0 U380 ( .INP(n148), .ZN(n323) );
  NOR2X0 U381 ( .IN1(n351), .IN2(n125), .QN(n195) );
  NOR2X0 U382 ( .IN1(n351), .IN2(instPacket_i[104]), .QN(n197) );
  INVX0 U383 ( .INP(instPacket_i[103]), .ZN(n351) );
  INVX0 U384 ( .INP(instPacket_i[101]), .ZN(n353) );
  NAND2X1 U385 ( .IN1(n201), .IN2(instPacket_i[101]), .QN(n173) );
  INVX0 U386 ( .INP(instPacket_i[102]), .ZN(n352) );
  INVX0 U387 ( .INP(instPacket_i[106]), .ZN(n340) );
  NOR2X0 U388 ( .IN1(instPacket_i[108]), .IN2(instPacket_i[107]), .QN(n202) );
  NBUFFX2 U389 ( .INP(instPacketValid_i), .Z(decodedPacket0Valid_o) );
  INVX0 U390 ( .INP(instPacket_i[105]), .ZN(n341) );
  INVX0 U391 ( .INP(instPacket_i[108]), .ZN(n328) );
  NOR4X0 U392 ( .IN1(n186), .IN2(instPacket_i[127]), .IN3(instPacket_i[129]), 
        .IN4(instPacket_i[128]), .QN(n185) );
  NOR4X0 U393 ( .IN1(n187), .IN2(instPacket_i[121]), .IN3(instPacket_i[123]), 
        .IN4(instPacket_i[122]), .QN(n184) );
  NOR4X0 U394 ( .IN1(n188), .IN2(instPacket_i[115]), .IN3(instPacket_i[117]), 
        .IN4(instPacket_i[116]), .QN(n183) );
  NOR4X0 U395 ( .IN1(n189), .IN2(instPacket_i[109]), .IN3(instPacket_i[111]), 
        .IN4(instPacket_i[110]), .QN(n182) );
  NOR4X0 U396 ( .IN1(n92), .IN2(n91), .IN3(n306), .IN4(n123), .QN(n122) );
  INVX0 U397 ( .INP(n128), .ZN(n346) );
  NOR2X0 U398 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[102]), .QN(n127) );
  NOR2X0 U399 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[103]), .QN(n128) );
  NAND2X1 U400 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[104]), .QN(n125)
         );
  NOR2X0 U401 ( .IN1(n125), .IN2(instPacket_i[101]), .QN(n131) );
  INVX0 U402 ( .INP(instPacket_i[107]), .ZN(n339) );
  INVX0 U403 ( .INP(instPacket_i_90), .ZN(n356) );
  NAND2X1 U404 ( .IN1(n324), .IN2(instPacket_i[101]), .QN(n148) );
  NBUFFX2 U405 ( .INP(instPacket_i[38]), .Z(decodedPacket0_o[38]) );
  NBUFFX2 U406 ( .INP(instPacket_i[39]), .Z(decodedPacket0_o[39]) );
  NBUFFX2 U407 ( .INP(instPacket_i[40]), .Z(decodedPacket0_o[40]) );
  NBUFFX2 U408 ( .INP(instPacket_i[41]), .Z(decodedPacket0_o[41]) );
  NBUFFX2 U409 ( .INP(instPacket_i[42]), .Z(decodedPacket0_o[42]) );
  NBUFFX2 U410 ( .INP(instPacket_i[43]), .Z(decodedPacket0_o[43]) );
  NBUFFX2 U411 ( .INP(instPacket_i[44]), .Z(decodedPacket0_o[44]) );
  NBUFFX2 U412 ( .INP(instPacket_i[45]), .Z(decodedPacket0_o[45]) );
  NBUFFX2 U413 ( .INP(instPacket_i[46]), .Z(decodedPacket0_o[46]) );
  NBUFFX2 U414 ( .INP(instPacket_i[47]), .Z(decodedPacket0_o[47]) );
  NBUFFX2 U415 ( .INP(instPacket_i[48]), .Z(decodedPacket0_o[48]) );
  NBUFFX2 U416 ( .INP(instPacket_i[49]), .Z(decodedPacket0_o[49]) );
  NBUFFX2 U417 ( .INP(instPacket_i[50]), .Z(decodedPacket0_o[50]) );
  NBUFFX2 U418 ( .INP(instPacket_i[51]), .Z(decodedPacket0_o[51]) );
  NBUFFX2 U419 ( .INP(instPacket_i[52]), .Z(decodedPacket0_o[52]) );
  NBUFFX2 U420 ( .INP(instPacket_i[53]), .Z(decodedPacket0_o[53]) );
  NBUFFX2 U421 ( .INP(instPacket_i[54]), .Z(decodedPacket0_o[54]) );
  NBUFFX2 U422 ( .INP(instPacket_i[55]), .Z(decodedPacket0_o[55]) );
  NBUFFX2 U423 ( .INP(instPacket_i[56]), .Z(decodedPacket0_o[56]) );
  NBUFFX2 U424 ( .INP(instPacket_i[57]), .Z(decodedPacket0_o[57]) );
  NBUFFX2 U425 ( .INP(instPacket_i[58]), .Z(decodedPacket0_o[58]) );
  NBUFFX2 U426 ( .INP(instPacket_i[59]), .Z(decodedPacket0_o[59]) );
  NBUFFX2 U427 ( .INP(instPacket_i[60]), .Z(decodedPacket0_o[60]) );
  NBUFFX2 U428 ( .INP(instPacket_i[61]), .Z(decodedPacket0_o[61]) );
  NBUFFX2 U429 ( .INP(instPacket_i[62]), .Z(decodedPacket0_o[62]) );
  NBUFFX2 U430 ( .INP(instPacket_i[63]), .Z(decodedPacket0_o[63]) );
  NBUFFX2 U431 ( .INP(instPacket_i[64]), .Z(decodedPacket0_o[64]) );
  NBUFFX2 U432 ( .INP(instPacket_i[65]), .Z(decodedPacket0_o[65]) );
  NBUFFX2 U433 ( .INP(instPacket_i[66]), .Z(decodedPacket0_o[66]) );
  NBUFFX2 U434 ( .INP(instPacket_i[67]), .Z(decodedPacket0_o[67]) );
  NBUFFX2 U435 ( .INP(instPacket_i[68]), .Z(decodedPacket0_o[68]) );
  NOR2X0 U436 ( .IN1(n138), .IN2(n353), .QN(n137) );
  NBUFFX2 U437 ( .INP(instPacket_i[0]), .Z(decodedPacket0_o[0]) );
  NBUFFX2 U438 ( .INP(instPacket_i[1]), .Z(decodedPacket0_o[1]) );
  NBUFFX2 U439 ( .INP(instPacket_i[2]), .Z(decodedPacket0_o[2]) );
  NBUFFX2 U440 ( .INP(instPacket_i[3]), .Z(decodedPacket0_o[3]) );
  NBUFFX2 U441 ( .INP(instPacket_i[4]), .Z(decodedPacket0_o[4]) );
  NBUFFX2 U442 ( .INP(instPacket_i[37]), .Z(decodedPacket0_o[37]) );
  NOR4X0 U443 ( .IN1(n70), .IN2(n71), .IN3(n72), .IN4(n73), .QN(n68) );
  NOR2X0 U444 ( .IN1(n74), .IN2(n356), .QN(n71) );
  INVX0 U445 ( .INP(instPacket_i_85), .ZN(n361) );
  INVX0 U446 ( .INP(instPacket_i_93), .ZN(n355) );
  INVX0 U447 ( .INP(instPacket_i_98), .ZN(n354) );
  INVX0 U448 ( .INP(instPacket_i_77), .ZN(n369) );
  INVX0 U449 ( .INP(instPacket_i_78), .ZN(n368) );
  INVX0 U450 ( .INP(instPacket_i_79), .ZN(n367) );
  INVX0 U451 ( .INP(instPacket_i_80), .ZN(n366) );
  INVX0 U452 ( .INP(instPacket_i_81), .ZN(n365) );
  INVX0 U453 ( .INP(instPacket_i_86), .ZN(n360) );
  INVX0 U454 ( .INP(instPacket_i_87), .ZN(n359) );
  INVX0 U455 ( .INP(instPacket_i_88), .ZN(n358) );
  INVX0 U456 ( .INP(instPacket_i_89), .ZN(n357) );
  INVX0 U457 ( .INP(instPacket_i_71), .ZN(N287) );
  INVX0 U458 ( .INP(instPacket_i_82), .ZN(n364) );
  INVX0 U459 ( .INP(instPacket_i_83), .ZN(n363) );
  INVX0 U460 ( .INP(instPacket_i_84), .ZN(n362) );
  NBUFFX2 U461 ( .INP(instPacket_i[1]), .Z(decodedPacket1_o[1]) );
  NBUFFX2 U462 ( .INP(instPacket_i[2]), .Z(decodedPacket1_o[2]) );
  NBUFFX2 U463 ( .INP(instPacket_i[3]), .Z(decodedPacket1_o[3]) );
  NBUFFX2 U464 ( .INP(instPacket_i[4]), .Z(decodedPacket1_o[4]) );
  NBUFFX2 U465 ( .INP(instPacket_i[37]), .Z(decodedPacket1_o[37]) );
  NBUFFX2 U466 ( .INP(instPacket_i[38]), .Z(decodedPacket1_o[38]) );
  NBUFFX2 U467 ( .INP(instPacket_i[39]), .Z(decodedPacket1_o[39]) );
  NBUFFX2 U468 ( .INP(instPacket_i[40]), .Z(decodedPacket1_o[40]) );
  NBUFFX2 U469 ( .INP(instPacket_i[41]), .Z(decodedPacket1_o[41]) );
  NBUFFX2 U470 ( .INP(instPacket_i[42]), .Z(decodedPacket1_o[42]) );
  NBUFFX2 U471 ( .INP(instPacket_i[43]), .Z(decodedPacket1_o[43]) );
  NBUFFX2 U472 ( .INP(instPacket_i[44]), .Z(decodedPacket1_o[44]) );
  NBUFFX2 U473 ( .INP(instPacket_i[45]), .Z(decodedPacket1_o[45]) );
  NBUFFX2 U474 ( .INP(instPacket_i[46]), .Z(decodedPacket1_o[46]) );
  NBUFFX2 U475 ( .INP(instPacket_i[47]), .Z(decodedPacket1_o[47]) );
  NBUFFX2 U476 ( .INP(instPacket_i[48]), .Z(decodedPacket1_o[48]) );
  NBUFFX2 U477 ( .INP(instPacket_i[49]), .Z(decodedPacket1_o[49]) );
  NBUFFX2 U478 ( .INP(instPacket_i[50]), .Z(decodedPacket1_o[50]) );
  NBUFFX2 U479 ( .INP(instPacket_i[51]), .Z(decodedPacket1_o[51]) );
  NBUFFX2 U480 ( .INP(instPacket_i[52]), .Z(decodedPacket1_o[52]) );
  NBUFFX2 U481 ( .INP(instPacket_i[53]), .Z(decodedPacket1_o[53]) );
  NBUFFX2 U482 ( .INP(instPacket_i[54]), .Z(decodedPacket1_o[54]) );
  NBUFFX2 U483 ( .INP(instPacket_i[55]), .Z(decodedPacket1_o[55]) );
  NBUFFX2 U484 ( .INP(instPacket_i[56]), .Z(decodedPacket1_o[56]) );
  NBUFFX2 U485 ( .INP(instPacket_i[57]), .Z(decodedPacket1_o[57]) );
  NBUFFX2 U486 ( .INP(instPacket_i[58]), .Z(decodedPacket1_o[58]) );
  NBUFFX2 U487 ( .INP(instPacket_i[59]), .Z(decodedPacket1_o[59]) );
  NBUFFX2 U488 ( .INP(instPacket_i[60]), .Z(decodedPacket1_o[60]) );
  NBUFFX2 U489 ( .INP(instPacket_i[61]), .Z(decodedPacket1_o[61]) );
  NBUFFX2 U490 ( .INP(instPacket_i[62]), .Z(decodedPacket1_o[62]) );
  NBUFFX2 U491 ( .INP(instPacket_i[63]), .Z(decodedPacket1_o[63]) );
  NBUFFX2 U492 ( .INP(instPacket_i[64]), .Z(decodedPacket1_o[64]) );
  NBUFFX2 U493 ( .INP(instPacket_i[65]), .Z(decodedPacket1_o[65]) );
  NBUFFX2 U494 ( .INP(instPacket_i[66]), .Z(decodedPacket1_o[66]) );
  NBUFFX2 U495 ( .INP(instPacket_i[67]), .Z(decodedPacket1_o[67]) );
  NBUFFX2 U496 ( .INP(instPacket_i[68]), .Z(decodedPacket1_o[68]) );
  NBUFFX2 U497 ( .INP(instPacket_i[0]), .Z(decodedPacket1_o[0]) );
  NBUFFX2 U498 ( .INP(n67), .Z(n311) );
  NBUFFX2 U499 ( .INP(n370), .Z(decodedPacket0_o[121]) );
  NAND4X0 U500 ( .IN1(n182), .IN2(n183), .IN3(n184), .IN4(n185), .QN(n306) );
  NAND4X0 U501 ( .IN1(n182), .IN2(n183), .IN3(n184), .IN4(n185), .QN(n307) );
  XOR2X1 U502 ( .IN1(\r340/carry[15] ), .IN2(instPacket_i_84), .Q(N300) );
  AND2X1 U503 ( .IN1(instPacket_i_83), .IN2(\r340/carry[14] ), .Q(
        \r340/carry[15] ) );
  XOR2X1 U504 ( .IN1(\r340/carry[14] ), .IN2(instPacket_i_83), .Q(N299) );
  AND2X1 U505 ( .IN1(instPacket_i_82), .IN2(\r340/carry[13] ), .Q(
        \r340/carry[14] ) );
  XOR2X1 U506 ( .IN1(\r340/carry[13] ), .IN2(instPacket_i_82), .Q(N298) );
  AND2X1 U507 ( .IN1(instPacket_i_81), .IN2(\r340/carry[12] ), .Q(
        \r340/carry[13] ) );
  XOR2X1 U508 ( .IN1(\r340/carry[12] ), .IN2(instPacket_i_81), .Q(N297) );
  AND2X1 U509 ( .IN1(instPacket_i_80), .IN2(\r340/carry[11] ), .Q(
        \r340/carry[12] ) );
  XOR2X1 U510 ( .IN1(\r340/carry[11] ), .IN2(instPacket_i_80), .Q(N296) );
  AND2X1 U511 ( .IN1(instPacket_i_79), .IN2(\r340/carry[10] ), .Q(
        \r340/carry[11] ) );
  XOR2X1 U512 ( .IN1(\r340/carry[10] ), .IN2(instPacket_i_79), .Q(N295) );
  AND2X1 U513 ( .IN1(instPacket_i_78), .IN2(\r340/carry[9] ), .Q(
        \r340/carry[10] ) );
  XOR2X1 U514 ( .IN1(\r340/carry[9] ), .IN2(instPacket_i_78), .Q(N294) );
  AND2X1 U515 ( .IN1(instPacket_i_77), .IN2(\r340/carry[8] ), .Q(
        \r340/carry[9] ) );
  XOR2X1 U516 ( .IN1(\r340/carry[8] ), .IN2(instPacket_i_77), .Q(N293) );
  AND2X1 U517 ( .IN1(instPacket_i_76), .IN2(\r340/carry[7] ), .Q(
        \r340/carry[8] ) );
  XOR2X1 U518 ( .IN1(\r340/carry[7] ), .IN2(instPacket_i_76), .Q(N292) );
  AND2X1 U519 ( .IN1(instPacket_i_75), .IN2(\r340/carry[6] ), .Q(
        \r340/carry[7] ) );
  XOR2X1 U520 ( .IN1(\r340/carry[6] ), .IN2(instPacket_i_75), .Q(N291) );
  AND2X1 U521 ( .IN1(instPacket_i_74), .IN2(\r340/carry[5] ), .Q(
        \r340/carry[6] ) );
  XOR2X1 U522 ( .IN1(\r340/carry[5] ), .IN2(instPacket_i_74), .Q(N290) );
  AND2X1 U523 ( .IN1(instPacket_i_73), .IN2(\r340/carry[4] ), .Q(
        \r340/carry[5] ) );
  XOR2X1 U524 ( .IN1(\r340/carry[4] ), .IN2(instPacket_i_73), .Q(N289) );
  AND2X1 U525 ( .IN1(instPacket_i_72), .IN2(instPacket_i_71), .Q(
        \r340/carry[4] ) );
  XOR2X1 U526 ( .IN1(instPacket_i_71), .IN2(instPacket_i_72), .Q(N288) );
  XOR2X1 U527 ( .IN1(\r339/carry[5] ), .IN2(instPacket_i_90), .Q(N284) );
endmodule


module Decode_PISA_3 ( instPacketValid_i, instPacket_i, decodedPacket0Valid_o, 
        decodedPacket0_o, decodedPacket1Valid_o, decodedPacket1_o );
  input [132:0] instPacket_i;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  input instPacketValid_i;
  output decodedPacket0Valid_o, decodedPacket1Valid_o;
  wire   instPacket_i_98, instPacket_i_97, instPacket_i_96, instPacket_i_95,
         instPacket_i_94, instPacket_i_93, instPacket_i_92, instPacket_i_91,
         instPacket_i_90, instPacket_i_89, instPacket_i_88, instPacket_i_87,
         instPacket_i_86, instPacket_i_85, instPacket_i_84, instPacket_i_83,
         instPacket_i_82, instPacket_i_81, instPacket_i_80, instPacket_i_79,
         instPacket_i_78, instPacket_i_77, instPacket_i_76, instPacket_i_75,
         instPacket_i_74, instPacket_i_73, instPacket_i_72, instPacket_i_71,
         instPacket_i_36, instPacket_i_35, instPacket_i_34, instPacket_i_33,
         instPacket_i_32, instPacket_i_31, instPacket_i_30, instPacket_i_29,
         instPacket_i_28, instPacket_i_27, instPacket_i_26, instPacket_i_25,
         instPacket_i_24, instPacket_i_23, instPacket_i_22, instPacket_i_21,
         instPacket_i_20, instPacket_i_19, instPacket_i_18, instPacket_i_17,
         instPacket_i_16, instPacket_i_15, instPacket_i_14, instPacket_i_13,
         instPacket_i_12, instPacket_i_11, instPacket_i_10, instPacket_i_9,
         instPacket_i_8, instPacket_i_7, instPacket_i_6, instPacket_i_5, n510,
         decodedPacket1_o_120, decodedPacket1_o_119, decodedPacket1_o_118,
         n511, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         \r340/carry[14] , \r340/carry[13] , \r340/carry[12] ,
         \r340/carry[11] , \r340/carry[10] , \r340/carry[9] , \r340/carry[8] ,
         \r340/carry[7] , \r340/carry[6] , \r340/carry[5] , \r340/carry[4] ,
         \r339/carry[5] , \r339/carry[4] , \r339/carry[3] , \r339/carry[2] ,
         n224, n225, n307, n308, n312, n313, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509;
  assign instPacket_i_98 = instPacket_i[98];
  assign instPacket_i_97 = instPacket_i[97];
  assign instPacket_i_96 = instPacket_i[96];
  assign instPacket_i_95 = instPacket_i[95];
  assign instPacket_i_94 = instPacket_i[94];
  assign instPacket_i_93 = instPacket_i[93];
  assign instPacket_i_92 = instPacket_i[92];
  assign instPacket_i_91 = instPacket_i[91];
  assign instPacket_i_90 = instPacket_i[90];
  assign instPacket_i_89 = instPacket_i[89];
  assign instPacket_i_88 = instPacket_i[88];
  assign instPacket_i_87 = instPacket_i[87];
  assign instPacket_i_86 = instPacket_i[86];
  assign instPacket_i_85 = instPacket_i[85];
  assign instPacket_i_84 = instPacket_i[84];
  assign instPacket_i_83 = instPacket_i[83];
  assign instPacket_i_82 = instPacket_i[82];
  assign instPacket_i_81 = instPacket_i[81];
  assign instPacket_i_80 = instPacket_i[80];
  assign instPacket_i_79 = instPacket_i[79];
  assign instPacket_i_78 = instPacket_i[78];
  assign instPacket_i_77 = instPacket_i[77];
  assign instPacket_i_76 = instPacket_i[76];
  assign instPacket_i_75 = instPacket_i[75];
  assign instPacket_i_74 = instPacket_i[74];
  assign instPacket_i_73 = instPacket_i[73];
  assign instPacket_i_72 = instPacket_i[72];
  assign instPacket_i_71 = instPacket_i[71];
  assign instPacket_i_36 = instPacket_i[36];
  assign instPacket_i_35 = instPacket_i[35];
  assign instPacket_i_34 = instPacket_i[34];
  assign instPacket_i_33 = instPacket_i[33];
  assign instPacket_i_32 = instPacket_i[32];
  assign instPacket_i_31 = instPacket_i[31];
  assign instPacket_i_30 = instPacket_i[30];
  assign instPacket_i_29 = instPacket_i[29];
  assign instPacket_i_28 = instPacket_i[28];
  assign instPacket_i_27 = instPacket_i[27];
  assign instPacket_i_26 = instPacket_i[26];
  assign instPacket_i_25 = instPacket_i[25];
  assign instPacket_i_24 = instPacket_i[24];
  assign instPacket_i_23 = instPacket_i[23];
  assign instPacket_i_22 = instPacket_i[22];
  assign instPacket_i_21 = instPacket_i[21];
  assign instPacket_i_20 = instPacket_i[20];
  assign instPacket_i_19 = instPacket_i[19];
  assign instPacket_i_18 = instPacket_i[18];
  assign instPacket_i_17 = instPacket_i[17];
  assign instPacket_i_16 = instPacket_i[16];
  assign instPacket_i_15 = instPacket_i[15];
  assign instPacket_i_14 = instPacket_i[14];
  assign instPacket_i_13 = instPacket_i[13];
  assign instPacket_i_12 = instPacket_i[12];
  assign instPacket_i_11 = instPacket_i[11];
  assign instPacket_i_10 = instPacket_i[10];
  assign instPacket_i_9 = instPacket_i[9];
  assign instPacket_i_8 = instPacket_i[8];
  assign instPacket_i_7 = instPacket_i[7];
  assign instPacket_i_6 = instPacket_i[6];
  assign instPacket_i_5 = instPacket_i[5];
  assign decodedPacket1_o[120] = decodedPacket1_o_120;
  assign decodedPacket1_o[119] = decodedPacket1_o_119;
  assign decodedPacket1_o[116] = decodedPacket1_o_118;
  assign N285 = instPacket_i[69];
  assign N286 = instPacket_i[70];

  AND2X1 U160 ( .IN1(N285), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[99]) );
  AO21X1 U161 ( .IN1(N284), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[97]) );
  AND2X1 U162 ( .IN1(decodedPacket1_o_119), .IN2(N283), .Q(
        decodedPacket1_o[96]) );
  AND2X1 U163 ( .IN1(decodedPacket1_o_119), .IN2(N282), .Q(
        decodedPacket1_o[95]) );
  AND2X1 U164 ( .IN1(decodedPacket1_o_119), .IN2(N281), .Q(
        decodedPacket1_o[94]) );
  AND2X1 U165 ( .IN1(decodedPacket1_o_119), .IN2(N280), .Q(
        decodedPacket1_o[93]) );
  AO21X1 U166 ( .IN1(n362), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[92]) );
  OR2X1 U167 ( .IN1(decodedPacket1_o_119), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[91]) );
  AO22X1 U168 ( .IN1(decodedPacket1_o_120), .IN2(N284), .IN3(instPacket_i_90), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[90]) );
  AO22X1 U169 ( .IN1(decodedPacket1_o_120), .IN2(N283), .IN3(instPacket_i_89), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[89]) );
  AO22X1 U170 ( .IN1(decodedPacket1_o_120), .IN2(N282), .IN3(instPacket_i_88), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[88]) );
  AO22X1 U171 ( .IN1(decodedPacket1_o_120), .IN2(N281), .IN3(instPacket_i_87), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[87]) );
  AO22X1 U172 ( .IN1(decodedPacket1_o_120), .IN2(N280), .IN3(instPacket_i_86), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[86]) );
  AO22X1 U173 ( .IN1(decodedPacket1_o_120), .IN2(n362), .IN3(instPacket_i_85), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[85]) );
  OR2X1 U174 ( .IN1(decodedPacket1_o_120), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[84]) );
  AND2X1 U175 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_97), .Q(
        decodedPacket1_o[82]) );
  AND2X1 U176 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_96), .Q(
        decodedPacket1_o[81]) );
  AND2X1 U177 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_95), .Q(
        decodedPacket1_o[80]) );
  AND2X1 U178 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_94), .Q(
        decodedPacket1_o[79]) );
  AND2X1 U179 ( .IN1(N300), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[114]) );
  AND2X1 U180 ( .IN1(N299), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[113]) );
  AND2X1 U181 ( .IN1(N298), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[112]) );
  AND2X1 U182 ( .IN1(N297), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[111]) );
  AND2X1 U183 ( .IN1(N296), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[110]) );
  AND2X1 U184 ( .IN1(N295), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[109]) );
  AND2X1 U185 ( .IN1(N294), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[108]) );
  AND2X1 U186 ( .IN1(N293), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[107]) );
  AND2X1 U187 ( .IN1(N292), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[106]) );
  AND2X1 U188 ( .IN1(N291), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[105]) );
  AND2X1 U189 ( .IN1(N290), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[104]) );
  AND2X1 U190 ( .IN1(N289), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[103]) );
  AND2X1 U191 ( .IN1(N288), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[102]) );
  AND2X1 U192 ( .IN1(N287), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[101]) );
  AND2X1 U193 ( .IN1(N286), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[100]) );
  AND2X1 U194 ( .IN1(instPacketValid_i), .IN2(decodedPacket1_o[76]), .Q(
        decodedPacket1Valid_o) );
  AO22X1 U195 ( .IN1(instPacket_i_9), .IN2(n510), .IN3(instPacket_i_73), .IN4(
        n312), .Q(decodedPacket0_o[9]) );
  AND2X1 U196 ( .IN1(decodedPacket0_o[98]), .IN2(N285), .Q(
        decodedPacket0_o[99]) );
  AO21X1 U197 ( .IN1(instPacket_i_82), .IN2(n500), .IN3(n499), .Q(n505) );
  OA221X1 U198 ( .IN1(n318), .IN2(n366), .IN3(n501), .IN4(n358), .IN5(n339), 
        .Q(n498) );
  OA221X1 U199 ( .IN1(n318), .IN2(n367), .IN3(n501), .IN4(n359), .IN5(n339), 
        .Q(n497) );
  OA221X1 U200 ( .IN1(n318), .IN2(n368), .IN3(n501), .IN4(n360), .IN5(n339), 
        .Q(n496) );
  OA221X1 U201 ( .IN1(n318), .IN2(n369), .IN3(n501), .IN4(n361), .IN5(n339), 
        .Q(n495) );
  OA221X1 U202 ( .IN1(n318), .IN2(n370), .IN3(n501), .IN4(n362), .IN5(n493), 
        .Q(n494) );
  AND3X1 U203 ( .IN1(n491), .IN2(n336), .IN3(n334), .Q(n501) );
  NAND4X0 U204 ( .IN1(n490), .IN2(n319), .IN3(n489), .IN4(n488), .QN(n500) );
  NAND4X0 U205 ( .IN1(n489), .IN2(n339), .IN3(n326), .IN4(n336), .QN(n486) );
  AO22X1 U206 ( .IN1(instPacket_i_8), .IN2(n510), .IN3(instPacket_i_72), .IN4(
        n508), .Q(decodedPacket0_o[8]) );
  NAND4X0 U207 ( .IN1(n490), .IN2(n331), .IN3(n323), .IN4(n480), .QN(n481) );
  NOR3X0 U208 ( .IN1(n479), .IN2(n333), .IN3(n478), .QN(n480) );
  OA21X1 U209 ( .IN1(n345), .IN2(n346), .IN3(n337), .Q(n479) );
  AND3X1 U210 ( .IN1(n477), .IN2(n320), .IN3(n327), .Q(n490) );
  OA221X1 U211 ( .IN1(n317), .IN2(n355), .IN3(n357), .IN4(n474), .IN5(n473), 
        .Q(n475) );
  AO22X1 U212 ( .IN1(n472), .IN2(instPacket_i_97), .IN3(n471), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[82]) );
  AO22X1 U213 ( .IN1(n472), .IN2(instPacket_i_96), .IN3(n471), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[81]) );
  AO22X1 U214 ( .IN1(n472), .IN2(instPacket_i_95), .IN3(n471), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[80]) );
  AO22X1 U215 ( .IN1(instPacket_i_7), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_71), .IN4(n508), .Q(decodedPacket0_o[7]) );
  AO22X1 U216 ( .IN1(n472), .IN2(instPacket_i_94), .IN3(n471), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[79]) );
  OA221X1 U217 ( .IN1(n317), .IN2(n356), .IN3(n362), .IN4(n474), .IN5(n469), 
        .Q(n470) );
  OA21X1 U218 ( .IN1(n467), .IN2(n468), .IN3(n315), .Q(decodedPacket0_o[77])
         );
  NAND4X0 U219 ( .IN1(n466), .IN2(n327), .IN3(n323), .IN4(n465), .QN(n468) );
  NAND3X0 U220 ( .IN1(n461), .IN2(n488), .IN3(n460), .QN(n485) );
  AO21X1 U221 ( .IN1(instPacket_i[104]), .IN2(n458), .IN3(decodedPacket1_o[72]), .Q(decodedPacket0_o[72]) );
  NAND3X0 U222 ( .IN1(n456), .IN2(n461), .IN3(n455), .QN(n457) );
  AO21X1 U223 ( .IN1(instPacket_i[102]), .IN2(n458), .IN3(decodedPacket1_o[70]), .Q(decodedPacket0_o[70]) );
  AO21X1 U224 ( .IN1(n315), .IN2(n321), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket1_o[70]) );
  AO22X1 U225 ( .IN1(instPacket_i_6), .IN2(decodedPacket0_o[121]), .IN3(N286), 
        .IN4(n508), .Q(decodedPacket0_o[6]) );
  AND2X1 U226 ( .IN1(n458), .IN2(instPacket_i[101]), .Q(decodedPacket0_o[69])
         );
  NAND4X0 U227 ( .IN1(n488), .IN2(n329), .IN3(n454), .IN4(n453), .QN(n458) );
  AND2X1 U228 ( .IN1(instPacket_i[106]), .IN2(n451), .Q(n452) );
  NAND4X0 U229 ( .IN1(n347), .IN2(n340), .IN3(n450), .IN4(n449), .QN(n451) );
  OA22X1 U230 ( .IN1(instPacket_i[105]), .IN2(n352), .IN3(n448), .IN4(n342), 
        .Q(n449) );
  AO22X1 U231 ( .IN1(n476), .IN2(n446), .IN3(n445), .IN4(n444), .Q(n484) );
  NAND4X0 U232 ( .IN1(n442), .IN2(n441), .IN3(n440), .IN4(n439), .QN(n446) );
  NOR3X0 U233 ( .IN1(n438), .IN2(n348), .IN3(n349), .QN(n439) );
  OA21X1 U234 ( .IN1(instPacket_i[103]), .IN2(n450), .IN3(n436), .Q(n437) );
  NAND4X0 U235 ( .IN1(n466), .IN2(n319), .IN3(n435), .IN4(n334), .QN(n483) );
  AND2X1 U236 ( .IN1(n320), .IN2(n434), .Q(n435) );
  OA21X1 U237 ( .IN1(n348), .IN2(n349), .IN3(n325), .Q(n463) );
  AND2X1 U238 ( .IN1(n469), .IN2(n433), .Q(n473) );
  NAND3X0 U239 ( .IN1(n325), .IN2(n354), .IN3(n351), .QN(n433) );
  OR2X1 U240 ( .IN1(n440), .IN2(n443), .Q(n469) );
  AND4X1 U241 ( .IN1(n432), .IN2(n431), .IN3(n430), .IN4(n429), .Q(n466) );
  NOR3X0 U242 ( .IN1(n450), .IN2(instPacket_i[103]), .IN3(n427), .QN(n503) );
  AOI22X1 U243 ( .IN1(n340), .IN2(n341), .IN3(instPacket_i[103]), .IN4(
        instPacket_i[104]), .QN(n454) );
  OR2X1 U244 ( .IN1(n443), .IN2(n426), .Q(n488) );
  AO22X1 U245 ( .IN1(instPacket_i_5), .IN2(n510), .IN3(N285), .IN4(n508), .Q(
        decodedPacket0_o[5]) );
  AND2X1 U246 ( .IN1(instPacket_i_36), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[36]) );
  AND2X1 U247 ( .IN1(instPacket_i_35), .IN2(n510), .Q(decodedPacket0_o[35]) );
  AND2X1 U248 ( .IN1(instPacket_i_34), .IN2(n510), .Q(decodedPacket0_o[34]) );
  AND2X1 U249 ( .IN1(instPacket_i_33), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[33]) );
  AND2X1 U250 ( .IN1(instPacket_i_32), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[32]) );
  AND2X1 U251 ( .IN1(instPacket_i_31), .IN2(n510), .Q(decodedPacket0_o[31]) );
  AO22X1 U252 ( .IN1(instPacket_i_30), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_94), .Q(decodedPacket0_o[30]) );
  AO22X1 U253 ( .IN1(instPacket_i_29), .IN2(n313), .IN3(n508), .IN4(
        instPacket_i_93), .Q(decodedPacket0_o[29]) );
  AO22X1 U254 ( .IN1(instPacket_i_28), .IN2(n313), .IN3(instPacket_i_92), 
        .IN4(n508), .Q(decodedPacket0_o[28]) );
  AO22X1 U255 ( .IN1(instPacket_i_27), .IN2(n313), .IN3(instPacket_i_91), 
        .IN4(n508), .Q(decodedPacket0_o[27]) );
  AO22X1 U256 ( .IN1(instPacket_i_26), .IN2(n313), .IN3(n508), .IN4(
        instPacket_i_90), .Q(decodedPacket0_o[26]) );
  AO22X1 U257 ( .IN1(instPacket_i_25), .IN2(n313), .IN3(n312), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[25]) );
  AO22X1 U258 ( .IN1(instPacket_i_24), .IN2(n313), .IN3(n508), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[24]) );
  AO22X1 U259 ( .IN1(instPacket_i_23), .IN2(n313), .IN3(n312), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[23]) );
  AO22X1 U260 ( .IN1(instPacket_i_22), .IN2(n313), .IN3(n508), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[22]) );
  AO22X1 U261 ( .IN1(instPacket_i_21), .IN2(n313), .IN3(n508), .IN4(
        instPacket_i_85), .Q(decodedPacket0_o[21]) );
  AO22X1 U262 ( .IN1(instPacket_i_20), .IN2(n313), .IN3(instPacket_i_84), 
        .IN4(n312), .Q(decodedPacket0_o[20]) );
  AO22X1 U263 ( .IN1(instPacket_i_19), .IN2(n313), .IN3(instPacket_i_83), 
        .IN4(n312), .Q(decodedPacket0_o[19]) );
  AO22X1 U264 ( .IN1(instPacket_i_18), .IN2(n313), .IN3(instPacket_i_82), 
        .IN4(n312), .Q(decodedPacket0_o[18]) );
  AO22X1 U265 ( .IN1(instPacket_i_17), .IN2(n313), .IN3(instPacket_i_81), 
        .IN4(n312), .Q(decodedPacket0_o[17]) );
  AO22X1 U266 ( .IN1(instPacket_i_16), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_80), .IN4(n312), .Q(decodedPacket0_o[16]) );
  AO22X1 U267 ( .IN1(instPacket_i_15), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_79), .IN4(n312), .Q(decodedPacket0_o[15]) );
  AO22X1 U268 ( .IN1(instPacket_i_14), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_78), .IN4(n312), .Q(decodedPacket0_o[14]) );
  AO22X1 U269 ( .IN1(instPacket_i_13), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_77), .IN4(n312), .Q(decodedPacket0_o[13]) );
  AO22X1 U270 ( .IN1(instPacket_i_12), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_76), .IN4(n312), .Q(decodedPacket0_o[12]) );
  AO21X1 U271 ( .IN1(n315), .IN2(n425), .IN3(decodedPacket1_o_120), .Q(
        decodedPacket0_o[120]) );
  AO22X1 U272 ( .IN1(instPacket_i_11), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_75), .IN4(n312), .Q(decodedPacket0_o[11]) );
  AO21X1 U273 ( .IN1(n315), .IN2(n423), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket0_o[119]) );
  NOR3X0 U275 ( .IN1(n419), .IN2(n332), .IN3(n418), .QN(n420) );
  NAND3X0 U276 ( .IN1(n413), .IN2(n338), .IN3(n455), .QN(n415) );
  NAND3X0 U277 ( .IN1(n426), .IN2(n410), .IN3(n409), .QN(n411) );
  AND2X1 U278 ( .IN1(n315), .IN2(n408), .Q(decodedPacket0_o[115]) );
  NAND4X0 U279 ( .IN1(n459), .IN2(n334), .IN3(n331), .IN4(n407), .QN(n408) );
  NAND4X0 U280 ( .IN1(n349), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n407) );
  AND2X1 U281 ( .IN1(n455), .IN2(n322), .Q(n459) );
  NAND3X0 U282 ( .IN1(n326), .IN2(n461), .IN3(n460), .QN(n499) );
  OA21X1 U283 ( .IN1(n441), .IN2(n443), .IN3(n456), .Q(n460) );
  OR2X1 U284 ( .IN1(n443), .IN2(n404), .Q(n461) );
  AO22X1 U285 ( .IN1(instPacket_i_10), .IN2(n313), .IN3(instPacket_i_74), 
        .IN4(n312), .Q(decodedPacket0_o[10]) );
  AND2X1 U286 ( .IN1(n315), .IN2(n414), .Q(n508) );
  AO21X1 U287 ( .IN1(n337), .IN2(n401), .IN3(n492), .Q(n414) );
  OA21X1 U288 ( .IN1(n464), .IN2(n412), .IN3(n315), .Q(n510) );
  AND2X1 U289 ( .IN1(n337), .IN2(n398), .Q(n464) );
  NAND4X0 U290 ( .IN1(n426), .IN2(n428), .IN3(n397), .IN4(n404), .QN(n398) );
  AND2X1 U291 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_76), .Q(
        decodedPacket0_o[106]) );
  AND2X1 U292 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_75), .Q(
        decodedPacket0_o[105]) );
  AND2X1 U293 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_74), .Q(
        decodedPacket0_o[104]) );
  AND2X1 U294 ( .IN1(instPacket_i_73), .IN2(decodedPacket0_o[98]), .Q(
        decodedPacket0_o[103]) );
  AND2X1 U295 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_72), .Q(
        decodedPacket0_o[102]) );
  AND2X1 U296 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_71), .Q(
        decodedPacket0_o[101]) );
  AND2X1 U297 ( .IN1(decodedPacket0_o[98]), .IN2(N286), .Q(
        decodedPacket0_o[100]) );
  NAND4X0 U299 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n506) );
  OR3X1 U300 ( .IN1(instPacket_i[132]), .IN2(instPacket_i[131]), .IN3(
        instPacket_i[130]), .Q(n390) );
  OR3X1 U301 ( .IN1(instPacket_i[126]), .IN2(instPacket_i[125]), .IN3(
        instPacket_i[124]), .Q(n389) );
  OR3X1 U302 ( .IN1(instPacket_i[120]), .IN2(instPacket_i[119]), .IN3(
        instPacket_i[118]), .Q(n388) );
  OR3X1 U303 ( .IN1(instPacket_i[114]), .IN2(instPacket_i[113]), .IN3(
        instPacket_i[112]), .Q(n387) );
  NAND3X0 U304 ( .IN1(n403), .IN2(n385), .IN3(n404), .QN(n386) );
  NAND3X0 U305 ( .IN1(n330), .IN2(n384), .IN3(n491), .QN(n395) );
  AND4X1 U306 ( .IN1(n432), .IN2(n431), .IN3(n383), .IN4(n434), .Q(n491) );
  NAND4X0 U307 ( .IN1(n348), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n434) );
  AOI22X1 U308 ( .IN1(n401), .IN2(n325), .IN3(n476), .IN4(n382), .QN(n431) );
  AO22X1 U309 ( .IN1(n351), .IN2(n354), .IN3(n444), .IN4(instPacket_i[103]), 
        .Q(n382) );
  NAND3X0 U310 ( .IN1(instPacket_i[103]), .IN2(n353), .IN3(instPacket_i[104]), 
        .QN(n436) );
  AOI222X1 U311 ( .IN1(n476), .IN2(n401), .IN3(n381), .IN4(n324), .IN5(n350), 
        .IN6(n325), .QN(n432) );
  NAND3X0 U312 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[101]), .IN3(n447), 
        .QN(n410) );
  AND3X1 U313 ( .IN1(instPacket_i[101]), .IN2(n353), .IN3(n447), .Q(n401) );
  AND2X1 U314 ( .IN1(n380), .IN2(instPacket_i[105]), .Q(n476) );
  AND3X1 U315 ( .IN1(n341), .IN2(n329), .IN3(instPacket_i[107]), .Q(n380) );
  AO21X1 U316 ( .IN1(n409), .IN2(n385), .IN3(n399), .Q(n384) );
  AND3X1 U317 ( .IN1(n396), .IN2(n404), .IN3(n397), .Q(n409) );
  AND2X1 U318 ( .IN1(n441), .IN2(n403), .Q(n397) );
  NAND3X0 U319 ( .IN1(instPacket_i[101]), .IN2(n379), .IN3(instPacket_i[102]), 
        .QN(n404) );
  NAND4X0 U320 ( .IN1(n331), .IN2(n406), .IN3(n378), .IN4(n455), .QN(n462) );
  NAND3X0 U321 ( .IN1(n379), .IN2(n353), .IN3(instPacket_i[101]), .QN(n385) );
  AND3X1 U322 ( .IN1(n353), .IN2(n352), .IN3(instPacket_i[104]), .Q(n375) );
  NAND3X0 U323 ( .IN1(n342), .IN2(n341), .IN3(n374), .QN(n399) );
  NOR3X0 U324 ( .IN1(n419), .IN2(n418), .IN3(n373), .QN(n406) );
  AOI21X1 U325 ( .IN1(n400), .IN2(n372), .IN3(n376), .QN(n373) );
  NAND3X0 U326 ( .IN1(n374), .IN2(n342), .IN3(instPacket_i[106]), .QN(n376) );
  NAND3X0 U327 ( .IN1(n379), .IN2(n354), .IN3(instPacket_i[102]), .QN(n396) );
  NAND3X0 U328 ( .IN1(n421), .IN2(n417), .IN3(n371), .QN(n425) );
  NAND3X0 U329 ( .IN1(n354), .IN2(n353), .IN3(n447), .QN(n372) );
  NAND3X0 U330 ( .IN1(instPacket_i[102]), .IN2(n354), .IN3(n447), .QN(n400) );
  AND3X1 U331 ( .IN1(instPacket_i[105]), .IN2(n374), .IN3(instPacket_i[106]), 
        .Q(n377) );
  NAND3X0 U332 ( .IN1(n354), .IN2(n353), .IN3(n379), .QN(n442) );
  HADDX1 \r339/U1_1_1  ( .A0(instPacket_i_86), .B0(instPacket_i_85), .C1(
        \r339/carry[2] ), .SO(N280) );
  HADDX1 \r339/U1_1_2  ( .A0(instPacket_i_87), .B0(\r339/carry[2] ), .C1(
        \r339/carry[3] ), .SO(N281) );
  HADDX1 \r339/U1_1_3  ( .A0(instPacket_i_88), .B0(\r339/carry[3] ), .C1(
        \r339/carry[4] ), .SO(N282) );
  HADDX1 \r339/U1_1_4  ( .A0(instPacket_i_89), .B0(\r339/carry[4] ), .C1(
        \r339/carry[5] ), .SO(N283) );
  INVX0 U3 ( .INP(1'b1), .ZN(decodedPacket1_o[5]) );
  INVX0 U5 ( .INP(1'b1), .ZN(decodedPacket1_o[6]) );
  INVX0 U7 ( .INP(1'b1), .ZN(decodedPacket1_o[7]) );
  INVX0 U9 ( .INP(1'b1), .ZN(decodedPacket1_o[8]) );
  INVX0 U11 ( .INP(1'b1), .ZN(decodedPacket1_o[9]) );
  INVX0 U13 ( .INP(1'b1), .ZN(decodedPacket1_o[10]) );
  INVX0 U15 ( .INP(1'b1), .ZN(decodedPacket1_o[11]) );
  INVX0 U17 ( .INP(1'b1), .ZN(decodedPacket1_o[12]) );
  INVX0 U19 ( .INP(1'b1), .ZN(decodedPacket1_o[13]) );
  INVX0 U21 ( .INP(1'b1), .ZN(decodedPacket1_o[14]) );
  INVX0 U23 ( .INP(1'b1), .ZN(decodedPacket1_o[15]) );
  INVX0 U25 ( .INP(1'b1), .ZN(decodedPacket1_o[16]) );
  INVX0 U27 ( .INP(1'b1), .ZN(decodedPacket1_o[17]) );
  INVX0 U29 ( .INP(1'b1), .ZN(decodedPacket1_o[18]) );
  INVX0 U31 ( .INP(1'b1), .ZN(decodedPacket1_o[19]) );
  INVX0 U33 ( .INP(1'b1), .ZN(decodedPacket1_o[20]) );
  INVX0 U35 ( .INP(1'b1), .ZN(decodedPacket1_o[21]) );
  INVX0 U37 ( .INP(1'b1), .ZN(decodedPacket1_o[22]) );
  INVX0 U39 ( .INP(1'b1), .ZN(decodedPacket1_o[23]) );
  INVX0 U41 ( .INP(1'b1), .ZN(decodedPacket1_o[24]) );
  INVX0 U43 ( .INP(1'b1), .ZN(decodedPacket1_o[25]) );
  INVX0 U45 ( .INP(1'b1), .ZN(decodedPacket1_o[26]) );
  INVX0 U47 ( .INP(1'b1), .ZN(decodedPacket1_o[27]) );
  INVX0 U49 ( .INP(1'b1), .ZN(decodedPacket1_o[28]) );
  INVX0 U51 ( .INP(1'b1), .ZN(decodedPacket1_o[29]) );
  INVX0 U53 ( .INP(1'b1), .ZN(decodedPacket1_o[30]) );
  INVX0 U55 ( .INP(1'b1), .ZN(decodedPacket1_o[31]) );
  INVX0 U57 ( .INP(1'b1), .ZN(decodedPacket1_o[32]) );
  INVX0 U59 ( .INP(1'b1), .ZN(decodedPacket1_o[33]) );
  INVX0 U61 ( .INP(1'b1), .ZN(decodedPacket1_o[34]) );
  INVX0 U63 ( .INP(1'b1), .ZN(decodedPacket1_o[35]) );
  INVX0 U65 ( .INP(1'b1), .ZN(decodedPacket1_o[36]) );
  INVX0 U67 ( .INP(1'b1), .ZN(decodedPacket1_o[117]) );
  INVX0 U69 ( .INP(1'b1), .ZN(decodedPacket1_o[121]) );
  INVX0 U71 ( .INP(1'b1), .ZN(decodedPacket1_o[122]) );
  INVX0 U73 ( .INP(1'b1), .ZN(decodedPacket1_o[123]) );
  INVX0 U75 ( .INP(1'b1), .ZN(decodedPacket1_o[124]) );
  INVX0 U77 ( .INP(1'b1), .ZN(decodedPacket1_o[125]) );
  INVX0 U79 ( .INP(1'b1), .ZN(decodedPacket0_o[122]) );
  INVX0 U81 ( .INP(1'b1), .ZN(decodedPacket0_o[123]) );
  INVX0 U83 ( .INP(1'b1), .ZN(decodedPacket0_o[124]) );
  INVX0 U85 ( .INP(1'b1), .ZN(decodedPacket0_o[125]) );
  INVX0 U87 ( .INP(decodedPacket1_o[77]), .ZN(n316) );
  NBUFFX2 U88 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[73]) );
  NBUFFX2 U89 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[75]) );
  NBUFFX2 U90 ( .INP(decodedPacket1_o[76]), .Z(decodedPacket1_o[115]) );
  NBUFFX2 U91 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[69]) );
  NBUFFX2 U92 ( .INP(n511), .Z(decodedPacket1_o[76]) );
  NBUFFX2 U93 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[98]) );
  NBUFFX2 U94 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[118]) );
  NBUFFX2 U95 ( .INP(n511), .Z(decodedPacket1_o[74]) );
  NBUFFX2 U96 ( .INP(n511), .Z(decodedPacket1_o[77]) );
  NOR2X0 U97 ( .IN1(n506), .IN2(n459), .QN(n511) );
  INVX0 U98 ( .INP(n499), .ZN(n322) );
  NOR2X0 U99 ( .IN1(n336), .IN2(n308), .QN(decodedPacket1_o_119) );
  INVX0 U100 ( .INP(n509), .ZN(decodedPacket1_o[71]) );
  NBUFFX2 U101 ( .INP(n510), .Z(decodedPacket0_o[121]) );
  INVX0 U102 ( .INP(n468), .ZN(n317) );
  INVX0 U103 ( .INP(n500), .ZN(n318) );
  NOR2X0 U104 ( .IN1(n308), .IN2(n317), .QN(n472) );
  INVX0 U105 ( .INP(n482), .ZN(decodedPacket0_o[84]) );
  INVX0 U106 ( .INP(n460), .ZN(n321) );
  NAND2X1 U107 ( .IN1(n343), .IN2(n337), .QN(n489) );
  INVX0 U108 ( .INP(n423), .ZN(n334) );
  INVX0 U109 ( .INP(n485), .ZN(n323) );
  INVX0 U110 ( .INP(n467), .ZN(n319) );
  INVX0 U111 ( .INP(n463), .ZN(n320) );
  NOR2X0 U112 ( .IN1(n422), .IN2(n333), .QN(n455) );
  INVX0 U113 ( .INP(n424), .ZN(n333) );
  NAND2X1 U114 ( .IN1(n345), .IN2(n325), .QN(n456) );
  INVX0 U115 ( .INP(n478), .ZN(n326) );
  INVX0 U116 ( .INP(n443), .ZN(n325) );
  NOR2X0 U117 ( .IN1(n307), .IN2(n322), .QN(decodedPacket1_o[72]) );
  NOR2X0 U118 ( .IN1(n308), .IN2(n455), .QN(decodedPacket1_o_118) );
  NAND2X1 U119 ( .IN1(n315), .IN2(n395), .QN(n402) );
  NAND2X1 U120 ( .IN1(n315), .IN2(n481), .QN(n482) );
  INVX0 U121 ( .INP(n506), .ZN(n315) );
  NOR2X0 U122 ( .IN1(n412), .IN2(n405), .QN(n378) );
  NOR4X0 U123 ( .IN1(n464), .IN2(n463), .IN3(n478), .IN4(n462), .QN(n465) );
  NOR2X0 U124 ( .IN1(n307), .IN2(n424), .QN(decodedPacket1_o_120) );
  INVX0 U125 ( .INP(n399), .ZN(n337) );
  INVX0 U126 ( .INP(n442), .ZN(n343) );
  NOR2X0 U127 ( .IN1(n440), .IN2(n399), .QN(n412) );
  NOR2X0 U128 ( .IN1(n420), .IN2(n307), .QN(decodedPacket0_o[117]) );
  INVX0 U129 ( .INP(n417), .ZN(n332) );
  INVX0 U130 ( .INP(n372), .ZN(n349) );
  INVX0 U131 ( .INP(n422), .ZN(n336) );
  NOR2X0 U132 ( .IN1(n474), .IN2(n308), .QN(n471) );
  NOR2X0 U133 ( .IN1(n343), .IN2(n346), .QN(n426) );
  OA21X1 U134 ( .IN1(n395), .IN2(n328), .IN3(n315), .Q(decodedPacket0_o[98])
         );
  INVX0 U135 ( .INP(n474), .ZN(n328) );
  NAND2X1 U136 ( .IN1(n406), .IN2(n335), .QN(n423) );
  INVX0 U137 ( .INP(n405), .ZN(n335) );
  INVX0 U138 ( .INP(n492), .ZN(n339) );
  NAND2X1 U139 ( .IN1(n315), .IN2(n457), .QN(n509) );
  NOR2X0 U140 ( .IN1(n350), .IN2(n345), .QN(n428) );
  INVX0 U141 ( .INP(n425), .ZN(n331) );
  NOR2X0 U142 ( .IN1(n416), .IN2(n307), .QN(decodedPacket0_o[116]) );
  NOR4X0 U143 ( .IN1(n415), .IN2(n414), .IN3(n425), .IN4(n423), .QN(n416) );
  INVX0 U144 ( .INP(n412), .ZN(n338) );
  NOR2X0 U145 ( .IN1(n487), .IN2(n307), .QN(decodedPacket0_o[91]) );
  NOR4X0 U146 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(n487) );
  NAND2X1 U147 ( .IN1(n473), .IN2(n474), .QN(n467) );
  OR2X1 U148 ( .IN1(decodedPacket1_o[118]), .IN2(n224), .Q(
        decodedPacket0_o[118]) );
  AOI21X1 U149 ( .IN1(n335), .IN2(n421), .IN3(n308), .QN(n224) );
  INVX0 U150 ( .INP(n484), .ZN(n327) );
  INVX0 U151 ( .INP(n396), .ZN(n345) );
  NOR2X0 U152 ( .IN1(n403), .IN2(n376), .QN(n422) );
  INVX0 U153 ( .INP(n385), .ZN(n346) );
  NOR2X0 U154 ( .IN1(n443), .IN2(n403), .QN(n478) );
  NAND2X1 U155 ( .IN1(n346), .IN2(n377), .QN(n424) );
  NAND2X1 U156 ( .IN1(n380), .IN2(n342), .QN(n443) );
  NAND2X1 U157 ( .IN1(n375), .IN2(n354), .QN(n441) );
  INVX0 U158 ( .INP(n462), .ZN(n330) );
  NAND2X1 U159 ( .IN1(n349), .IN2(n377), .QN(n371) );
  NOR2X0 U274 ( .IN1(n441), .IN2(n376), .QN(n405) );
  NOR2X0 U298 ( .IN1(n442), .IN2(n376), .QN(n418) );
  NOR2X0 U333 ( .IN1(n396), .IN2(n376), .QN(n419) );
  NOR2X0 U334 ( .IN1(n400), .IN2(n399), .QN(n492) );
  NAND2X1 U335 ( .IN1(n476), .IN2(n386), .QN(n474) );
  NOR2X0 U336 ( .IN1(n316), .IN2(n356), .QN(decodedPacket1_o[78]) );
  NOR2X0 U337 ( .IN1(n316), .IN2(n355), .QN(decodedPacket1_o[83]) );
  INVX0 U338 ( .INP(n400), .ZN(n348) );
  NOR2X0 U339 ( .IN1(n436), .IN2(n427), .QN(n502) );
  INVX0 U340 ( .INP(n410), .ZN(n350) );
  NOR2X0 U341 ( .IN1(n370), .IN2(n402), .QN(decodedPacket0_o[107]) );
  NOR2X0 U342 ( .IN1(n369), .IN2(n402), .QN(decodedPacket0_o[108]) );
  NOR2X0 U343 ( .IN1(n368), .IN2(n402), .QN(decodedPacket0_o[109]) );
  NOR2X0 U344 ( .IN1(n367), .IN2(n402), .QN(decodedPacket0_o[110]) );
  NOR2X0 U345 ( .IN1(n366), .IN2(n402), .QN(decodedPacket0_o[111]) );
  NOR2X0 U346 ( .IN1(n352), .IN2(n443), .QN(n445) );
  NOR2X0 U347 ( .IN1(n362), .IN2(n482), .QN(decodedPacket0_o[85]) );
  NOR2X0 U348 ( .IN1(n361), .IN2(n482), .QN(decodedPacket0_o[86]) );
  NOR2X0 U349 ( .IN1(n360), .IN2(n482), .QN(decodedPacket0_o[87]) );
  NOR2X0 U350 ( .IN1(n359), .IN2(n482), .QN(decodedPacket0_o[88]) );
  NOR2X0 U351 ( .IN1(n358), .IN2(n482), .QN(decodedPacket0_o[89]) );
  NOR2X0 U352 ( .IN1(n357), .IN2(n482), .QN(decodedPacket0_o[90]) );
  NAND2X1 U353 ( .IN1(n444), .IN2(n352), .QN(n440) );
  NAND2X1 U354 ( .IN1(n348), .IN2(n377), .QN(n417) );
  NOR2X0 U355 ( .IN1(n494), .IN2(n308), .QN(decodedPacket0_o[92]) );
  NOR2X0 U356 ( .IN1(n492), .IN2(n503), .QN(n493) );
  NOR2X0 U357 ( .IN1(n495), .IN2(n308), .QN(decodedPacket0_o[93]) );
  NOR2X0 U358 ( .IN1(n496), .IN2(n308), .QN(decodedPacket0_o[94]) );
  NOR2X0 U359 ( .IN1(n497), .IN2(n307), .QN(decodedPacket0_o[95]) );
  NOR2X0 U360 ( .IN1(n498), .IN2(n307), .QN(decodedPacket0_o[96]) );
  NOR2X0 U361 ( .IN1(n470), .IN2(n308), .QN(decodedPacket0_o[78]) );
  NOR2X0 U362 ( .IN1(n475), .IN2(n308), .QN(decodedPacket0_o[83]) );
  NAND2X1 U363 ( .IN1(n343), .IN2(n377), .QN(n421) );
  NAND2X1 U364 ( .IN1(n476), .IN2(n344), .QN(n429) );
  NOR2X0 U365 ( .IN1(n503), .IN2(n502), .QN(n430) );
  INVX0 U366 ( .INP(n428), .ZN(n344) );
  NAND2X1 U367 ( .IN1(n316), .IN2(n342), .QN(decodedPacket0_o[73]) );
  NAND2X1 U368 ( .IN1(n316), .IN2(n341), .QN(decodedPacket0_o[74]) );
  NAND2X1 U369 ( .IN1(n316), .IN2(n340), .QN(decodedPacket0_o[75]) );
  NAND2X1 U370 ( .IN1(n316), .IN2(n329), .QN(decodedPacket0_o[76]) );
  NAND2X1 U371 ( .IN1(n350), .IN2(n476), .QN(n383) );
  NAND2X1 U372 ( .IN1(n509), .IN2(n352), .QN(decodedPacket0_o[71]) );
  NAND2X1 U373 ( .IN1(n476), .IN2(n345), .QN(n477) );
  INVX0 U374 ( .INP(n436), .ZN(n351) );
  NAND2X1 U375 ( .IN1(n337), .IN2(n411), .QN(n413) );
  INVX0 U376 ( .INP(n427), .ZN(n324) );
  NOR2X0 U377 ( .IN1(n352), .IN2(n450), .QN(n381) );
  NOR2X0 U378 ( .IN1(n352), .IN2(instPacket_i[104]), .QN(n379) );
  NAND2X1 U379 ( .IN1(n375), .IN2(instPacket_i[101]), .QN(n403) );
  NBUFFX2 U380 ( .INP(instPacketValid_i), .Z(decodedPacket0Valid_o) );
  INVX0 U381 ( .INP(instPacket_i[103]), .ZN(n352) );
  INVX0 U382 ( .INP(instPacket_i[101]), .ZN(n354) );
  INVX0 U383 ( .INP(instPacket_i[105]), .ZN(n342) );
  INVX0 U384 ( .INP(instPacket_i[102]), .ZN(n353) );
  INVX0 U385 ( .INP(instPacket_i[106]), .ZN(n341) );
  NOR2X0 U386 ( .IN1(instPacket_i[108]), .IN2(instPacket_i[107]), .QN(n374) );
  INVX0 U387 ( .INP(instPacket_i[108]), .ZN(n329) );
  NOR4X0 U388 ( .IN1(n390), .IN2(instPacket_i[127]), .IN3(instPacket_i[129]), 
        .IN4(instPacket_i[128]), .QN(n391) );
  NOR4X0 U389 ( .IN1(n389), .IN2(instPacket_i[121]), .IN3(instPacket_i[123]), 
        .IN4(instPacket_i[122]), .QN(n392) );
  NOR4X0 U390 ( .IN1(n387), .IN2(instPacket_i[109]), .IN3(instPacket_i[111]), 
        .IN4(instPacket_i[110]), .QN(n394) );
  NOR4X0 U391 ( .IN1(n388), .IN2(instPacket_i[115]), .IN3(instPacket_i[117]), 
        .IN4(instPacket_i[116]), .QN(n393) );
  NOR4X0 U392 ( .IN1(n483), .IN2(n484), .IN3(n307), .IN4(n452), .QN(n453) );
  INVX0 U393 ( .INP(n447), .ZN(n347) );
  NOR2X0 U394 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[102]), .QN(n448) );
  INVX0 U395 ( .INP(instPacket_i_71), .ZN(N287) );
  XNOR2X1 U396 ( .IN1(n225), .IN2(instPacket_i_84), .Q(N300) );
  NAND2X1 U397 ( .IN1(instPacket_i_83), .IN2(\r340/carry[14] ), .QN(n225) );
  NOR2X0 U398 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[103]), .QN(n447) );
  NBUFFX2 U399 ( .INP(instPacket_i[0]), .Z(decodedPacket1_o[0]) );
  NBUFFX2 U400 ( .INP(instPacket_i[1]), .Z(decodedPacket1_o[1]) );
  NBUFFX2 U401 ( .INP(instPacket_i[2]), .Z(decodedPacket1_o[2]) );
  NBUFFX2 U402 ( .INP(instPacket_i[3]), .Z(decodedPacket1_o[3]) );
  NBUFFX2 U403 ( .INP(instPacket_i[4]), .Z(decodedPacket1_o[4]) );
  NBUFFX2 U404 ( .INP(instPacket_i[37]), .Z(decodedPacket1_o[37]) );
  NBUFFX2 U405 ( .INP(instPacket_i[38]), .Z(decodedPacket1_o[38]) );
  NBUFFX2 U406 ( .INP(instPacket_i[39]), .Z(decodedPacket1_o[39]) );
  NBUFFX2 U407 ( .INP(instPacket_i[40]), .Z(decodedPacket1_o[40]) );
  NBUFFX2 U408 ( .INP(instPacket_i[41]), .Z(decodedPacket1_o[41]) );
  NBUFFX2 U409 ( .INP(instPacket_i[42]), .Z(decodedPacket1_o[42]) );
  NBUFFX2 U410 ( .INP(instPacket_i[43]), .Z(decodedPacket1_o[43]) );
  NBUFFX2 U411 ( .INP(instPacket_i[44]), .Z(decodedPacket1_o[44]) );
  NBUFFX2 U412 ( .INP(instPacket_i[45]), .Z(decodedPacket1_o[45]) );
  NBUFFX2 U413 ( .INP(instPacket_i[46]), .Z(decodedPacket1_o[46]) );
  NBUFFX2 U414 ( .INP(instPacket_i[47]), .Z(decodedPacket1_o[47]) );
  NBUFFX2 U415 ( .INP(instPacket_i[48]), .Z(decodedPacket1_o[48]) );
  NBUFFX2 U416 ( .INP(instPacket_i[49]), .Z(decodedPacket1_o[49]) );
  NBUFFX2 U417 ( .INP(instPacket_i[50]), .Z(decodedPacket1_o[50]) );
  NBUFFX2 U418 ( .INP(instPacket_i[51]), .Z(decodedPacket1_o[51]) );
  NBUFFX2 U419 ( .INP(instPacket_i[52]), .Z(decodedPacket1_o[52]) );
  NBUFFX2 U420 ( .INP(instPacket_i[53]), .Z(decodedPacket1_o[53]) );
  NBUFFX2 U421 ( .INP(instPacket_i[54]), .Z(decodedPacket1_o[54]) );
  NBUFFX2 U422 ( .INP(instPacket_i[55]), .Z(decodedPacket1_o[55]) );
  NBUFFX2 U423 ( .INP(instPacket_i[56]), .Z(decodedPacket1_o[56]) );
  NBUFFX2 U424 ( .INP(instPacket_i[57]), .Z(decodedPacket1_o[57]) );
  NBUFFX2 U425 ( .INP(instPacket_i[58]), .Z(decodedPacket1_o[58]) );
  NBUFFX2 U426 ( .INP(instPacket_i[59]), .Z(decodedPacket1_o[59]) );
  NBUFFX2 U427 ( .INP(instPacket_i[60]), .Z(decodedPacket1_o[60]) );
  NBUFFX2 U428 ( .INP(instPacket_i[61]), .Z(decodedPacket1_o[61]) );
  NBUFFX2 U429 ( .INP(instPacket_i[62]), .Z(decodedPacket1_o[62]) );
  NBUFFX2 U430 ( .INP(instPacket_i[63]), .Z(decodedPacket1_o[63]) );
  NBUFFX2 U431 ( .INP(instPacket_i[64]), .Z(decodedPacket1_o[64]) );
  NBUFFX2 U432 ( .INP(instPacket_i[65]), .Z(decodedPacket1_o[65]) );
  NBUFFX2 U433 ( .INP(instPacket_i[66]), .Z(decodedPacket1_o[66]) );
  NBUFFX2 U434 ( .INP(instPacket_i[67]), .Z(decodedPacket1_o[67]) );
  NBUFFX2 U435 ( .INP(instPacket_i[68]), .Z(decodedPacket1_o[68]) );
  NOR2X0 U436 ( .IN1(n365), .IN2(n402), .QN(decodedPacket0_o[112]) );
  INVX0 U437 ( .INP(instPacket_i_82), .ZN(n365) );
  NOR2X0 U438 ( .IN1(n364), .IN2(n402), .QN(decodedPacket0_o[113]) );
  INVX0 U439 ( .INP(instPacket_i_83), .ZN(n364) );
  NOR2X0 U440 ( .IN1(n363), .IN2(n402), .QN(decodedPacket0_o[114]) );
  INVX0 U441 ( .INP(instPacket_i_84), .ZN(n363) );
  NAND2X1 U442 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[104]), .QN(n450)
         );
  NOR2X0 U443 ( .IN1(n450), .IN2(instPacket_i[101]), .QN(n444) );
  INVX0 U444 ( .INP(instPacket_i[107]), .ZN(n340) );
  INVX0 U445 ( .INP(instPacket_i_90), .ZN(n357) );
  NAND2X1 U446 ( .IN1(n325), .IN2(instPacket_i[101]), .QN(n427) );
  NOR2X0 U447 ( .IN1(n437), .IN2(n354), .QN(n438) );
  NOR2X0 U448 ( .IN1(n507), .IN2(n307), .QN(decodedPacket0_o[97]) );
  NOR4X0 U449 ( .IN1(n505), .IN2(n504), .IN3(n503), .IN4(n502), .QN(n507) );
  NOR2X0 U450 ( .IN1(n501), .IN2(n357), .QN(n504) );
  INVX0 U451 ( .INP(instPacket_i_85), .ZN(n362) );
  INVX0 U452 ( .INP(instPacket_i_93), .ZN(n356) );
  INVX0 U453 ( .INP(instPacket_i_98), .ZN(n355) );
  INVX0 U454 ( .INP(instPacket_i_77), .ZN(n370) );
  INVX0 U455 ( .INP(instPacket_i_78), .ZN(n369) );
  INVX0 U456 ( .INP(instPacket_i_79), .ZN(n368) );
  INVX0 U457 ( .INP(instPacket_i_80), .ZN(n367) );
  INVX0 U458 ( .INP(instPacket_i_81), .ZN(n366) );
  INVX0 U459 ( .INP(instPacket_i_86), .ZN(n361) );
  INVX0 U460 ( .INP(instPacket_i_87), .ZN(n360) );
  INVX0 U461 ( .INP(instPacket_i_88), .ZN(n359) );
  INVX0 U462 ( .INP(instPacket_i_89), .ZN(n358) );
  NBUFFX2 U463 ( .INP(instPacket_i[0]), .Z(decodedPacket0_o[0]) );
  NBUFFX2 U464 ( .INP(instPacket_i[1]), .Z(decodedPacket0_o[1]) );
  NBUFFX2 U465 ( .INP(instPacket_i[2]), .Z(decodedPacket0_o[2]) );
  NBUFFX2 U466 ( .INP(instPacket_i[3]), .Z(decodedPacket0_o[3]) );
  NBUFFX2 U467 ( .INP(instPacket_i[4]), .Z(decodedPacket0_o[4]) );
  NBUFFX2 U468 ( .INP(instPacket_i[37]), .Z(decodedPacket0_o[37]) );
  NBUFFX2 U469 ( .INP(instPacket_i[38]), .Z(decodedPacket0_o[38]) );
  NBUFFX2 U470 ( .INP(instPacket_i[39]), .Z(decodedPacket0_o[39]) );
  NBUFFX2 U471 ( .INP(instPacket_i[40]), .Z(decodedPacket0_o[40]) );
  NBUFFX2 U472 ( .INP(instPacket_i[41]), .Z(decodedPacket0_o[41]) );
  NBUFFX2 U473 ( .INP(instPacket_i[42]), .Z(decodedPacket0_o[42]) );
  NBUFFX2 U474 ( .INP(instPacket_i[43]), .Z(decodedPacket0_o[43]) );
  NBUFFX2 U475 ( .INP(instPacket_i[44]), .Z(decodedPacket0_o[44]) );
  NBUFFX2 U476 ( .INP(instPacket_i[45]), .Z(decodedPacket0_o[45]) );
  NBUFFX2 U477 ( .INP(instPacket_i[46]), .Z(decodedPacket0_o[46]) );
  NBUFFX2 U478 ( .INP(instPacket_i[47]), .Z(decodedPacket0_o[47]) );
  NBUFFX2 U479 ( .INP(instPacket_i[48]), .Z(decodedPacket0_o[48]) );
  NBUFFX2 U480 ( .INP(instPacket_i[49]), .Z(decodedPacket0_o[49]) );
  NBUFFX2 U481 ( .INP(instPacket_i[50]), .Z(decodedPacket0_o[50]) );
  NBUFFX2 U482 ( .INP(instPacket_i[51]), .Z(decodedPacket0_o[51]) );
  NBUFFX2 U483 ( .INP(instPacket_i[52]), .Z(decodedPacket0_o[52]) );
  NBUFFX2 U484 ( .INP(instPacket_i[53]), .Z(decodedPacket0_o[53]) );
  NBUFFX2 U485 ( .INP(instPacket_i[54]), .Z(decodedPacket0_o[54]) );
  NBUFFX2 U486 ( .INP(instPacket_i[55]), .Z(decodedPacket0_o[55]) );
  NBUFFX2 U487 ( .INP(instPacket_i[56]), .Z(decodedPacket0_o[56]) );
  NBUFFX2 U488 ( .INP(instPacket_i[57]), .Z(decodedPacket0_o[57]) );
  NBUFFX2 U489 ( .INP(instPacket_i[58]), .Z(decodedPacket0_o[58]) );
  NBUFFX2 U490 ( .INP(instPacket_i[59]), .Z(decodedPacket0_o[59]) );
  NBUFFX2 U491 ( .INP(instPacket_i[60]), .Z(decodedPacket0_o[60]) );
  NBUFFX2 U492 ( .INP(instPacket_i[61]), .Z(decodedPacket0_o[61]) );
  NBUFFX2 U493 ( .INP(instPacket_i[62]), .Z(decodedPacket0_o[62]) );
  NBUFFX2 U494 ( .INP(instPacket_i[63]), .Z(decodedPacket0_o[63]) );
  NBUFFX2 U495 ( .INP(instPacket_i[64]), .Z(decodedPacket0_o[64]) );
  NBUFFX2 U496 ( .INP(instPacket_i[65]), .Z(decodedPacket0_o[65]) );
  NBUFFX2 U497 ( .INP(instPacket_i[66]), .Z(decodedPacket0_o[66]) );
  NBUFFX2 U498 ( .INP(instPacket_i[67]), .Z(decodedPacket0_o[67]) );
  NBUFFX2 U499 ( .INP(instPacket_i[68]), .Z(decodedPacket0_o[68]) );
  NBUFFX2 U500 ( .INP(n508), .Z(n312) );
  NBUFFX2 U501 ( .INP(n510), .Z(n313) );
  NAND4X0 U502 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n307) );
  NAND4X0 U503 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n308) );
  XOR2X1 U504 ( .IN1(\r340/carry[14] ), .IN2(instPacket_i_83), .Q(N299) );
  AND2X1 U505 ( .IN1(instPacket_i_82), .IN2(\r340/carry[13] ), .Q(
        \r340/carry[14] ) );
  XOR2X1 U506 ( .IN1(\r340/carry[13] ), .IN2(instPacket_i_82), .Q(N298) );
  AND2X1 U507 ( .IN1(instPacket_i_81), .IN2(\r340/carry[12] ), .Q(
        \r340/carry[13] ) );
  XOR2X1 U508 ( .IN1(\r340/carry[12] ), .IN2(instPacket_i_81), .Q(N297) );
  AND2X1 U509 ( .IN1(instPacket_i_80), .IN2(\r340/carry[11] ), .Q(
        \r340/carry[12] ) );
  XOR2X1 U510 ( .IN1(\r340/carry[11] ), .IN2(instPacket_i_80), .Q(N296) );
  AND2X1 U511 ( .IN1(instPacket_i_79), .IN2(\r340/carry[10] ), .Q(
        \r340/carry[11] ) );
  XOR2X1 U512 ( .IN1(\r340/carry[10] ), .IN2(instPacket_i_79), .Q(N295) );
  AND2X1 U513 ( .IN1(instPacket_i_78), .IN2(\r340/carry[9] ), .Q(
        \r340/carry[10] ) );
  XOR2X1 U514 ( .IN1(\r340/carry[9] ), .IN2(instPacket_i_78), .Q(N294) );
  AND2X1 U515 ( .IN1(instPacket_i_77), .IN2(\r340/carry[8] ), .Q(
        \r340/carry[9] ) );
  XOR2X1 U516 ( .IN1(\r340/carry[8] ), .IN2(instPacket_i_77), .Q(N293) );
  AND2X1 U517 ( .IN1(instPacket_i_76), .IN2(\r340/carry[7] ), .Q(
        \r340/carry[8] ) );
  XOR2X1 U518 ( .IN1(\r340/carry[7] ), .IN2(instPacket_i_76), .Q(N292) );
  AND2X1 U519 ( .IN1(instPacket_i_75), .IN2(\r340/carry[6] ), .Q(
        \r340/carry[7] ) );
  XOR2X1 U520 ( .IN1(\r340/carry[6] ), .IN2(instPacket_i_75), .Q(N291) );
  AND2X1 U521 ( .IN1(instPacket_i_74), .IN2(\r340/carry[5] ), .Q(
        \r340/carry[6] ) );
  XOR2X1 U522 ( .IN1(\r340/carry[5] ), .IN2(instPacket_i_74), .Q(N290) );
  AND2X1 U523 ( .IN1(instPacket_i_73), .IN2(\r340/carry[4] ), .Q(
        \r340/carry[5] ) );
  XOR2X1 U524 ( .IN1(\r340/carry[4] ), .IN2(instPacket_i_73), .Q(N289) );
  AND2X1 U525 ( .IN1(instPacket_i_72), .IN2(instPacket_i_71), .Q(
        \r340/carry[4] ) );
  XOR2X1 U526 ( .IN1(instPacket_i_71), .IN2(instPacket_i_72), .Q(N288) );
  XOR2X1 U527 ( .IN1(\r339/carry[5] ), .IN2(instPacket_i_90), .Q(N284) );
endmodule


module Decode_PISA_2 ( instPacketValid_i, instPacket_i, decodedPacket0Valid_o, 
        decodedPacket0_o, decodedPacket1Valid_o, decodedPacket1_o );
  input [132:0] instPacket_i;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  input instPacketValid_i;
  output decodedPacket0Valid_o, decodedPacket1Valid_o;
  wire   instPacket_i_98, instPacket_i_97, instPacket_i_96, instPacket_i_95,
         instPacket_i_94, instPacket_i_93, instPacket_i_92, instPacket_i_91,
         instPacket_i_90, instPacket_i_89, instPacket_i_88, instPacket_i_87,
         instPacket_i_86, instPacket_i_85, instPacket_i_84, instPacket_i_83,
         instPacket_i_82, instPacket_i_81, instPacket_i_80, instPacket_i_79,
         instPacket_i_78, instPacket_i_77, instPacket_i_76, instPacket_i_75,
         instPacket_i_74, instPacket_i_73, instPacket_i_72, instPacket_i_71,
         instPacket_i_36, instPacket_i_35, instPacket_i_34, instPacket_i_33,
         instPacket_i_32, instPacket_i_31, instPacket_i_30, instPacket_i_29,
         instPacket_i_28, instPacket_i_27, instPacket_i_26, instPacket_i_25,
         instPacket_i_24, instPacket_i_23, instPacket_i_22, instPacket_i_21,
         instPacket_i_20, instPacket_i_19, instPacket_i_18, instPacket_i_17,
         instPacket_i_16, instPacket_i_15, instPacket_i_14, instPacket_i_13,
         instPacket_i_12, instPacket_i_11, instPacket_i_10, instPacket_i_9,
         instPacket_i_8, instPacket_i_7, instPacket_i_6, instPacket_i_5, n510,
         decodedPacket1_o_120, decodedPacket1_o_119, decodedPacket1_o_118,
         n511, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         \r340/carry[14] , \r340/carry[13] , \r340/carry[12] ,
         \r340/carry[11] , \r340/carry[10] , \r340/carry[9] , \r340/carry[8] ,
         \r340/carry[7] , \r340/carry[6] , \r340/carry[5] , \r340/carry[4] ,
         \r339/carry[5] , \r339/carry[4] , \r339/carry[3] , \r339/carry[2] ,
         n224, n225, n307, n308, n312, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509;
  assign instPacket_i_98 = instPacket_i[98];
  assign instPacket_i_97 = instPacket_i[97];
  assign instPacket_i_96 = instPacket_i[96];
  assign instPacket_i_95 = instPacket_i[95];
  assign instPacket_i_94 = instPacket_i[94];
  assign instPacket_i_93 = instPacket_i[93];
  assign instPacket_i_92 = instPacket_i[92];
  assign instPacket_i_91 = instPacket_i[91];
  assign instPacket_i_90 = instPacket_i[90];
  assign instPacket_i_89 = instPacket_i[89];
  assign instPacket_i_88 = instPacket_i[88];
  assign instPacket_i_87 = instPacket_i[87];
  assign instPacket_i_86 = instPacket_i[86];
  assign instPacket_i_85 = instPacket_i[85];
  assign instPacket_i_84 = instPacket_i[84];
  assign instPacket_i_83 = instPacket_i[83];
  assign instPacket_i_82 = instPacket_i[82];
  assign instPacket_i_81 = instPacket_i[81];
  assign instPacket_i_80 = instPacket_i[80];
  assign instPacket_i_79 = instPacket_i[79];
  assign instPacket_i_78 = instPacket_i[78];
  assign instPacket_i_77 = instPacket_i[77];
  assign instPacket_i_76 = instPacket_i[76];
  assign instPacket_i_75 = instPacket_i[75];
  assign instPacket_i_74 = instPacket_i[74];
  assign instPacket_i_73 = instPacket_i[73];
  assign instPacket_i_72 = instPacket_i[72];
  assign instPacket_i_71 = instPacket_i[71];
  assign instPacket_i_36 = instPacket_i[36];
  assign instPacket_i_35 = instPacket_i[35];
  assign instPacket_i_34 = instPacket_i[34];
  assign instPacket_i_33 = instPacket_i[33];
  assign instPacket_i_32 = instPacket_i[32];
  assign instPacket_i_31 = instPacket_i[31];
  assign instPacket_i_30 = instPacket_i[30];
  assign instPacket_i_29 = instPacket_i[29];
  assign instPacket_i_28 = instPacket_i[28];
  assign instPacket_i_27 = instPacket_i[27];
  assign instPacket_i_26 = instPacket_i[26];
  assign instPacket_i_25 = instPacket_i[25];
  assign instPacket_i_24 = instPacket_i[24];
  assign instPacket_i_23 = instPacket_i[23];
  assign instPacket_i_22 = instPacket_i[22];
  assign instPacket_i_21 = instPacket_i[21];
  assign instPacket_i_20 = instPacket_i[20];
  assign instPacket_i_19 = instPacket_i[19];
  assign instPacket_i_18 = instPacket_i[18];
  assign instPacket_i_17 = instPacket_i[17];
  assign instPacket_i_16 = instPacket_i[16];
  assign instPacket_i_15 = instPacket_i[15];
  assign instPacket_i_14 = instPacket_i[14];
  assign instPacket_i_13 = instPacket_i[13];
  assign instPacket_i_12 = instPacket_i[12];
  assign instPacket_i_11 = instPacket_i[11];
  assign instPacket_i_10 = instPacket_i[10];
  assign instPacket_i_9 = instPacket_i[9];
  assign instPacket_i_8 = instPacket_i[8];
  assign instPacket_i_7 = instPacket_i[7];
  assign instPacket_i_6 = instPacket_i[6];
  assign instPacket_i_5 = instPacket_i[5];
  assign decodedPacket1_o[120] = decodedPacket1_o_120;
  assign decodedPacket1_o[119] = decodedPacket1_o_119;
  assign decodedPacket1_o[116] = decodedPacket1_o_118;
  assign N285 = instPacket_i[69];
  assign N286 = instPacket_i[70];

  AND2X1 U160 ( .IN1(N285), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[99]) );
  AO21X1 U161 ( .IN1(N284), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[97]) );
  AND2X1 U162 ( .IN1(decodedPacket1_o_119), .IN2(N283), .Q(
        decodedPacket1_o[96]) );
  AND2X1 U163 ( .IN1(decodedPacket1_o_119), .IN2(N282), .Q(
        decodedPacket1_o[95]) );
  AND2X1 U164 ( .IN1(decodedPacket1_o_119), .IN2(N281), .Q(
        decodedPacket1_o[94]) );
  AND2X1 U165 ( .IN1(decodedPacket1_o_119), .IN2(N280), .Q(
        decodedPacket1_o[93]) );
  AO21X1 U166 ( .IN1(n362), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[92]) );
  OR2X1 U167 ( .IN1(decodedPacket1_o_119), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[91]) );
  AO22X1 U168 ( .IN1(decodedPacket1_o_120), .IN2(N284), .IN3(instPacket_i_90), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[90]) );
  AO22X1 U169 ( .IN1(decodedPacket1_o_120), .IN2(N283), .IN3(instPacket_i_89), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[89]) );
  AO22X1 U170 ( .IN1(decodedPacket1_o_120), .IN2(N282), .IN3(instPacket_i_88), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[88]) );
  AO22X1 U171 ( .IN1(decodedPacket1_o_120), .IN2(N281), .IN3(instPacket_i_87), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[87]) );
  AO22X1 U172 ( .IN1(decodedPacket1_o_120), .IN2(N280), .IN3(instPacket_i_86), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[86]) );
  AO22X1 U173 ( .IN1(decodedPacket1_o_120), .IN2(n362), .IN3(instPacket_i_85), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[85]) );
  OR2X1 U174 ( .IN1(decodedPacket1_o_120), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[84]) );
  AND2X1 U175 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_97), .Q(
        decodedPacket1_o[82]) );
  AND2X1 U176 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_96), .Q(
        decodedPacket1_o[81]) );
  AND2X1 U177 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_95), .Q(
        decodedPacket1_o[80]) );
  AND2X1 U178 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_94), .Q(
        decodedPacket1_o[79]) );
  AND2X1 U179 ( .IN1(N300), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[114]) );
  AND2X1 U180 ( .IN1(N299), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[113]) );
  AND2X1 U181 ( .IN1(N298), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[112]) );
  AND2X1 U182 ( .IN1(N297), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[111]) );
  AND2X1 U183 ( .IN1(N296), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[110]) );
  AND2X1 U184 ( .IN1(N295), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[109]) );
  AND2X1 U185 ( .IN1(N294), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[108]) );
  AND2X1 U186 ( .IN1(N293), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[107]) );
  AND2X1 U187 ( .IN1(N292), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[106]) );
  AND2X1 U188 ( .IN1(N291), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[105]) );
  AND2X1 U189 ( .IN1(N290), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[104]) );
  AND2X1 U190 ( .IN1(N289), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[103]) );
  AND2X1 U191 ( .IN1(N288), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[102]) );
  AND2X1 U192 ( .IN1(N287), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[101]) );
  AND2X1 U193 ( .IN1(N286), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[100]) );
  AND2X1 U194 ( .IN1(instPacketValid_i), .IN2(decodedPacket1_o[76]), .Q(
        decodedPacket1Valid_o) );
  AO22X1 U195 ( .IN1(instPacket_i_9), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_73), .IN4(n312), .Q(decodedPacket0_o[9]) );
  AND2X1 U196 ( .IN1(decodedPacket0_o[98]), .IN2(N285), .Q(
        decodedPacket0_o[99]) );
  AO21X1 U197 ( .IN1(instPacket_i_82), .IN2(n500), .IN3(n499), .Q(n505) );
  OA221X1 U198 ( .IN1(n318), .IN2(n366), .IN3(n501), .IN4(n358), .IN5(n339), 
        .Q(n498) );
  OA221X1 U199 ( .IN1(n318), .IN2(n367), .IN3(n501), .IN4(n359), .IN5(n339), 
        .Q(n497) );
  OA221X1 U200 ( .IN1(n318), .IN2(n368), .IN3(n501), .IN4(n360), .IN5(n339), 
        .Q(n496) );
  OA221X1 U201 ( .IN1(n318), .IN2(n369), .IN3(n501), .IN4(n361), .IN5(n339), 
        .Q(n495) );
  OA221X1 U202 ( .IN1(n318), .IN2(n370), .IN3(n501), .IN4(n362), .IN5(n493), 
        .Q(n494) );
  AND3X1 U203 ( .IN1(n491), .IN2(n336), .IN3(n334), .Q(n501) );
  NAND4X0 U204 ( .IN1(n490), .IN2(n319), .IN3(n489), .IN4(n488), .QN(n500) );
  NAND4X0 U205 ( .IN1(n489), .IN2(n339), .IN3(n326), .IN4(n336), .QN(n486) );
  AO22X1 U206 ( .IN1(instPacket_i_8), .IN2(n510), .IN3(instPacket_i_72), .IN4(
        n508), .Q(decodedPacket0_o[8]) );
  NAND4X0 U207 ( .IN1(n490), .IN2(n331), .IN3(n323), .IN4(n480), .QN(n481) );
  NOR3X0 U208 ( .IN1(n479), .IN2(n333), .IN3(n478), .QN(n480) );
  OA21X1 U209 ( .IN1(n345), .IN2(n346), .IN3(n337), .Q(n479) );
  AND3X1 U210 ( .IN1(n477), .IN2(n320), .IN3(n327), .Q(n490) );
  OA221X1 U211 ( .IN1(n317), .IN2(n355), .IN3(n357), .IN4(n474), .IN5(n473), 
        .Q(n475) );
  AO22X1 U212 ( .IN1(n472), .IN2(instPacket_i_97), .IN3(n471), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[82]) );
  AO22X1 U213 ( .IN1(n472), .IN2(instPacket_i_96), .IN3(n471), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[81]) );
  AO22X1 U214 ( .IN1(n472), .IN2(instPacket_i_95), .IN3(n471), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[80]) );
  AO22X1 U215 ( .IN1(instPacket_i_7), .IN2(n510), .IN3(instPacket_i_71), .IN4(
        n508), .Q(decodedPacket0_o[7]) );
  AO22X1 U216 ( .IN1(n472), .IN2(instPacket_i_94), .IN3(n471), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[79]) );
  OA221X1 U217 ( .IN1(n317), .IN2(n356), .IN3(n362), .IN4(n474), .IN5(n469), 
        .Q(n470) );
  OA21X1 U218 ( .IN1(n467), .IN2(n468), .IN3(n315), .Q(decodedPacket0_o[77])
         );
  NAND4X0 U219 ( .IN1(n466), .IN2(n327), .IN3(n323), .IN4(n465), .QN(n468) );
  NAND3X0 U220 ( .IN1(n461), .IN2(n488), .IN3(n460), .QN(n485) );
  AO21X1 U221 ( .IN1(instPacket_i[104]), .IN2(n458), .IN3(decodedPacket1_o[72]), .Q(decodedPacket0_o[72]) );
  NAND3X0 U222 ( .IN1(n456), .IN2(n461), .IN3(n455), .QN(n457) );
  AO21X1 U223 ( .IN1(instPacket_i[102]), .IN2(n458), .IN3(decodedPacket1_o[70]), .Q(decodedPacket0_o[70]) );
  AO21X1 U224 ( .IN1(n315), .IN2(n321), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket1_o[70]) );
  AO22X1 U225 ( .IN1(instPacket_i_6), .IN2(decodedPacket0_o[121]), .IN3(N286), 
        .IN4(n508), .Q(decodedPacket0_o[6]) );
  AND2X1 U226 ( .IN1(n458), .IN2(instPacket_i[101]), .Q(decodedPacket0_o[69])
         );
  NAND4X0 U227 ( .IN1(n488), .IN2(n329), .IN3(n454), .IN4(n453), .QN(n458) );
  AND2X1 U228 ( .IN1(instPacket_i[106]), .IN2(n451), .Q(n452) );
  NAND4X0 U229 ( .IN1(n347), .IN2(n340), .IN3(n450), .IN4(n449), .QN(n451) );
  OA22X1 U230 ( .IN1(instPacket_i[105]), .IN2(n352), .IN3(n448), .IN4(n342), 
        .Q(n449) );
  AO22X1 U231 ( .IN1(n476), .IN2(n446), .IN3(n445), .IN4(n444), .Q(n484) );
  NAND4X0 U232 ( .IN1(n442), .IN2(n441), .IN3(n440), .IN4(n439), .QN(n446) );
  NOR3X0 U233 ( .IN1(n438), .IN2(n348), .IN3(n349), .QN(n439) );
  OA21X1 U234 ( .IN1(instPacket_i[103]), .IN2(n450), .IN3(n436), .Q(n437) );
  NAND4X0 U235 ( .IN1(n466), .IN2(n319), .IN3(n435), .IN4(n334), .QN(n483) );
  AND2X1 U236 ( .IN1(n320), .IN2(n434), .Q(n435) );
  OA21X1 U237 ( .IN1(n348), .IN2(n349), .IN3(n325), .Q(n463) );
  AND2X1 U238 ( .IN1(n469), .IN2(n433), .Q(n473) );
  NAND3X0 U239 ( .IN1(n325), .IN2(n354), .IN3(n351), .QN(n433) );
  OR2X1 U240 ( .IN1(n440), .IN2(n443), .Q(n469) );
  AND4X1 U241 ( .IN1(n432), .IN2(n431), .IN3(n430), .IN4(n429), .Q(n466) );
  NOR3X0 U242 ( .IN1(n450), .IN2(instPacket_i[103]), .IN3(n427), .QN(n503) );
  AOI22X1 U243 ( .IN1(n340), .IN2(n341), .IN3(instPacket_i[103]), .IN4(
        instPacket_i[104]), .QN(n454) );
  OR2X1 U244 ( .IN1(n443), .IN2(n426), .Q(n488) );
  AO22X1 U245 ( .IN1(instPacket_i_5), .IN2(n510), .IN3(N285), .IN4(n508), .Q(
        decodedPacket0_o[5]) );
  AND2X1 U246 ( .IN1(instPacket_i_36), .IN2(n510), .Q(decodedPacket0_o[36]) );
  AND2X1 U247 ( .IN1(instPacket_i_35), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[35]) );
  AND2X1 U248 ( .IN1(instPacket_i_34), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[34]) );
  AND2X1 U249 ( .IN1(instPacket_i_33), .IN2(n510), .Q(decodedPacket0_o[33]) );
  AND2X1 U250 ( .IN1(instPacket_i_32), .IN2(n510), .Q(decodedPacket0_o[32]) );
  AND2X1 U251 ( .IN1(instPacket_i_31), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[31]) );
  AO22X1 U252 ( .IN1(instPacket_i_30), .IN2(n314), .IN3(n508), .IN4(
        instPacket_i_94), .Q(decodedPacket0_o[30]) );
  AO22X1 U253 ( .IN1(instPacket_i_29), .IN2(decodedPacket0_o[121]), .IN3(n508), 
        .IN4(instPacket_i_93), .Q(decodedPacket0_o[29]) );
  AO22X1 U254 ( .IN1(instPacket_i_28), .IN2(n510), .IN3(instPacket_i_92), 
        .IN4(n508), .Q(decodedPacket0_o[28]) );
  AO22X1 U255 ( .IN1(instPacket_i_27), .IN2(n314), .IN3(instPacket_i_91), 
        .IN4(n508), .Q(decodedPacket0_o[27]) );
  AO22X1 U256 ( .IN1(instPacket_i_26), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_90), .Q(decodedPacket0_o[26]) );
  AO22X1 U257 ( .IN1(instPacket_i_25), .IN2(n314), .IN3(n312), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[25]) );
  AO22X1 U258 ( .IN1(instPacket_i_24), .IN2(decodedPacket0_o[121]), .IN3(n508), 
        .IN4(instPacket_i_88), .Q(decodedPacket0_o[24]) );
  AO22X1 U259 ( .IN1(instPacket_i_23), .IN2(n510), .IN3(n312), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[23]) );
  AO22X1 U260 ( .IN1(instPacket_i_22), .IN2(n314), .IN3(n508), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[22]) );
  AO22X1 U261 ( .IN1(instPacket_i_21), .IN2(decodedPacket0_o[121]), .IN3(n508), 
        .IN4(instPacket_i_85), .Q(decodedPacket0_o[21]) );
  AO22X1 U262 ( .IN1(instPacket_i_20), .IN2(n314), .IN3(instPacket_i_84), 
        .IN4(n312), .Q(decodedPacket0_o[20]) );
  AO22X1 U263 ( .IN1(instPacket_i_19), .IN2(n314), .IN3(instPacket_i_83), 
        .IN4(n312), .Q(decodedPacket0_o[19]) );
  AO22X1 U264 ( .IN1(instPacket_i_18), .IN2(n314), .IN3(instPacket_i_82), 
        .IN4(n312), .Q(decodedPacket0_o[18]) );
  AO22X1 U265 ( .IN1(instPacket_i_17), .IN2(n314), .IN3(instPacket_i_81), 
        .IN4(n312), .Q(decodedPacket0_o[17]) );
  AO22X1 U266 ( .IN1(instPacket_i_16), .IN2(n314), .IN3(instPacket_i_80), 
        .IN4(n312), .Q(decodedPacket0_o[16]) );
  AO22X1 U267 ( .IN1(instPacket_i_15), .IN2(n314), .IN3(instPacket_i_79), 
        .IN4(n312), .Q(decodedPacket0_o[15]) );
  AO22X1 U268 ( .IN1(instPacket_i_14), .IN2(n314), .IN3(instPacket_i_78), 
        .IN4(n312), .Q(decodedPacket0_o[14]) );
  AO22X1 U269 ( .IN1(instPacket_i_13), .IN2(n314), .IN3(instPacket_i_77), 
        .IN4(n312), .Q(decodedPacket0_o[13]) );
  AO22X1 U270 ( .IN1(instPacket_i_12), .IN2(n314), .IN3(instPacket_i_76), 
        .IN4(n312), .Q(decodedPacket0_o[12]) );
  AO21X1 U271 ( .IN1(n315), .IN2(n425), .IN3(decodedPacket1_o_120), .Q(
        decodedPacket0_o[120]) );
  AO22X1 U272 ( .IN1(instPacket_i_11), .IN2(n314), .IN3(instPacket_i_75), 
        .IN4(n312), .Q(decodedPacket0_o[11]) );
  AO21X1 U273 ( .IN1(n315), .IN2(n423), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket0_o[119]) );
  NOR3X0 U275 ( .IN1(n419), .IN2(n332), .IN3(n418), .QN(n420) );
  NAND3X0 U276 ( .IN1(n413), .IN2(n338), .IN3(n455), .QN(n415) );
  NAND3X0 U277 ( .IN1(n426), .IN2(n410), .IN3(n409), .QN(n411) );
  AND2X1 U278 ( .IN1(n315), .IN2(n408), .Q(decodedPacket0_o[115]) );
  NAND4X0 U279 ( .IN1(n459), .IN2(n334), .IN3(n331), .IN4(n407), .QN(n408) );
  NAND4X0 U280 ( .IN1(n349), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n407) );
  AND2X1 U281 ( .IN1(n455), .IN2(n322), .Q(n459) );
  NAND3X0 U282 ( .IN1(n326), .IN2(n461), .IN3(n460), .QN(n499) );
  OA21X1 U283 ( .IN1(n441), .IN2(n443), .IN3(n456), .Q(n460) );
  OR2X1 U284 ( .IN1(n443), .IN2(n404), .Q(n461) );
  AO22X1 U285 ( .IN1(instPacket_i_10), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_74), .IN4(n312), .Q(decodedPacket0_o[10]) );
  AND2X1 U286 ( .IN1(n315), .IN2(n414), .Q(n508) );
  AO21X1 U287 ( .IN1(n337), .IN2(n401), .IN3(n492), .Q(n414) );
  OA21X1 U288 ( .IN1(n464), .IN2(n412), .IN3(n315), .Q(n510) );
  AND2X1 U289 ( .IN1(n337), .IN2(n398), .Q(n464) );
  NAND4X0 U290 ( .IN1(n426), .IN2(n428), .IN3(n397), .IN4(n404), .QN(n398) );
  AND2X1 U291 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_76), .Q(
        decodedPacket0_o[106]) );
  AND2X1 U292 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_75), .Q(
        decodedPacket0_o[105]) );
  AND2X1 U293 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_74), .Q(
        decodedPacket0_o[104]) );
  AND2X1 U294 ( .IN1(instPacket_i_73), .IN2(decodedPacket0_o[98]), .Q(
        decodedPacket0_o[103]) );
  AND2X1 U295 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_72), .Q(
        decodedPacket0_o[102]) );
  AND2X1 U296 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_71), .Q(
        decodedPacket0_o[101]) );
  AND2X1 U297 ( .IN1(decodedPacket0_o[98]), .IN2(N286), .Q(
        decodedPacket0_o[100]) );
  NAND4X0 U299 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n506) );
  OR3X1 U300 ( .IN1(instPacket_i[132]), .IN2(instPacket_i[131]), .IN3(
        instPacket_i[130]), .Q(n390) );
  OR3X1 U301 ( .IN1(instPacket_i[126]), .IN2(instPacket_i[125]), .IN3(
        instPacket_i[124]), .Q(n389) );
  OR3X1 U302 ( .IN1(instPacket_i[120]), .IN2(instPacket_i[119]), .IN3(
        instPacket_i[118]), .Q(n388) );
  OR3X1 U303 ( .IN1(instPacket_i[114]), .IN2(instPacket_i[113]), .IN3(
        instPacket_i[112]), .Q(n387) );
  NAND3X0 U304 ( .IN1(n403), .IN2(n385), .IN3(n404), .QN(n386) );
  NAND3X0 U305 ( .IN1(n330), .IN2(n384), .IN3(n491), .QN(n395) );
  AND4X1 U306 ( .IN1(n432), .IN2(n431), .IN3(n383), .IN4(n434), .Q(n491) );
  NAND4X0 U307 ( .IN1(n348), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n434) );
  AOI22X1 U308 ( .IN1(n401), .IN2(n325), .IN3(n476), .IN4(n382), .QN(n431) );
  AO22X1 U309 ( .IN1(n351), .IN2(n354), .IN3(n444), .IN4(instPacket_i[103]), 
        .Q(n382) );
  NAND3X0 U310 ( .IN1(instPacket_i[103]), .IN2(n353), .IN3(instPacket_i[104]), 
        .QN(n436) );
  AOI222X1 U311 ( .IN1(n476), .IN2(n401), .IN3(n381), .IN4(n324), .IN5(n350), 
        .IN6(n325), .QN(n432) );
  NAND3X0 U312 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[101]), .IN3(n447), 
        .QN(n410) );
  AND3X1 U313 ( .IN1(instPacket_i[101]), .IN2(n353), .IN3(n447), .Q(n401) );
  AND2X1 U314 ( .IN1(n380), .IN2(instPacket_i[105]), .Q(n476) );
  AND3X1 U315 ( .IN1(n341), .IN2(n329), .IN3(instPacket_i[107]), .Q(n380) );
  AO21X1 U316 ( .IN1(n409), .IN2(n385), .IN3(n399), .Q(n384) );
  AND3X1 U317 ( .IN1(n396), .IN2(n404), .IN3(n397), .Q(n409) );
  AND2X1 U318 ( .IN1(n441), .IN2(n403), .Q(n397) );
  NAND3X0 U319 ( .IN1(instPacket_i[101]), .IN2(n379), .IN3(instPacket_i[102]), 
        .QN(n404) );
  NAND4X0 U320 ( .IN1(n331), .IN2(n406), .IN3(n378), .IN4(n455), .QN(n462) );
  NAND3X0 U321 ( .IN1(n379), .IN2(n353), .IN3(instPacket_i[101]), .QN(n385) );
  AND3X1 U322 ( .IN1(n353), .IN2(n352), .IN3(instPacket_i[104]), .Q(n375) );
  NAND3X0 U323 ( .IN1(n342), .IN2(n341), .IN3(n374), .QN(n399) );
  NOR3X0 U324 ( .IN1(n419), .IN2(n418), .IN3(n373), .QN(n406) );
  AOI21X1 U325 ( .IN1(n400), .IN2(n372), .IN3(n376), .QN(n373) );
  NAND3X0 U326 ( .IN1(n374), .IN2(n342), .IN3(instPacket_i[106]), .QN(n376) );
  NAND3X0 U327 ( .IN1(n379), .IN2(n354), .IN3(instPacket_i[102]), .QN(n396) );
  NAND3X0 U328 ( .IN1(n421), .IN2(n417), .IN3(n371), .QN(n425) );
  NAND3X0 U329 ( .IN1(n354), .IN2(n353), .IN3(n447), .QN(n372) );
  NAND3X0 U330 ( .IN1(instPacket_i[102]), .IN2(n354), .IN3(n447), .QN(n400) );
  AND3X1 U331 ( .IN1(instPacket_i[105]), .IN2(n374), .IN3(instPacket_i[106]), 
        .Q(n377) );
  NAND3X0 U332 ( .IN1(n354), .IN2(n353), .IN3(n379), .QN(n442) );
  HADDX1 \r339/U1_1_1  ( .A0(instPacket_i_86), .B0(instPacket_i_85), .C1(
        \r339/carry[2] ), .SO(N280) );
  HADDX1 \r339/U1_1_2  ( .A0(instPacket_i_87), .B0(\r339/carry[2] ), .C1(
        \r339/carry[3] ), .SO(N281) );
  HADDX1 \r339/U1_1_3  ( .A0(instPacket_i_88), .B0(\r339/carry[3] ), .C1(
        \r339/carry[4] ), .SO(N282) );
  HADDX1 \r339/U1_1_4  ( .A0(instPacket_i_89), .B0(\r339/carry[4] ), .C1(
        \r339/carry[5] ), .SO(N283) );
  INVX0 U3 ( .INP(1'b1), .ZN(decodedPacket1_o[5]) );
  INVX0 U5 ( .INP(1'b1), .ZN(decodedPacket1_o[6]) );
  INVX0 U7 ( .INP(1'b1), .ZN(decodedPacket1_o[7]) );
  INVX0 U9 ( .INP(1'b1), .ZN(decodedPacket1_o[8]) );
  INVX0 U11 ( .INP(1'b1), .ZN(decodedPacket1_o[9]) );
  INVX0 U13 ( .INP(1'b1), .ZN(decodedPacket1_o[10]) );
  INVX0 U15 ( .INP(1'b1), .ZN(decodedPacket1_o[11]) );
  INVX0 U17 ( .INP(1'b1), .ZN(decodedPacket1_o[12]) );
  INVX0 U19 ( .INP(1'b1), .ZN(decodedPacket1_o[13]) );
  INVX0 U21 ( .INP(1'b1), .ZN(decodedPacket1_o[14]) );
  INVX0 U23 ( .INP(1'b1), .ZN(decodedPacket1_o[15]) );
  INVX0 U25 ( .INP(1'b1), .ZN(decodedPacket1_o[16]) );
  INVX0 U27 ( .INP(1'b1), .ZN(decodedPacket1_o[17]) );
  INVX0 U29 ( .INP(1'b1), .ZN(decodedPacket1_o[18]) );
  INVX0 U31 ( .INP(1'b1), .ZN(decodedPacket1_o[19]) );
  INVX0 U33 ( .INP(1'b1), .ZN(decodedPacket1_o[20]) );
  INVX0 U35 ( .INP(1'b1), .ZN(decodedPacket1_o[21]) );
  INVX0 U37 ( .INP(1'b1), .ZN(decodedPacket1_o[22]) );
  INVX0 U39 ( .INP(1'b1), .ZN(decodedPacket1_o[23]) );
  INVX0 U41 ( .INP(1'b1), .ZN(decodedPacket1_o[24]) );
  INVX0 U43 ( .INP(1'b1), .ZN(decodedPacket1_o[25]) );
  INVX0 U45 ( .INP(1'b1), .ZN(decodedPacket1_o[26]) );
  INVX0 U47 ( .INP(1'b1), .ZN(decodedPacket1_o[27]) );
  INVX0 U49 ( .INP(1'b1), .ZN(decodedPacket1_o[28]) );
  INVX0 U51 ( .INP(1'b1), .ZN(decodedPacket1_o[29]) );
  INVX0 U53 ( .INP(1'b1), .ZN(decodedPacket1_o[30]) );
  INVX0 U55 ( .INP(1'b1), .ZN(decodedPacket1_o[31]) );
  INVX0 U57 ( .INP(1'b1), .ZN(decodedPacket1_o[32]) );
  INVX0 U59 ( .INP(1'b1), .ZN(decodedPacket1_o[33]) );
  INVX0 U61 ( .INP(1'b1), .ZN(decodedPacket1_o[34]) );
  INVX0 U63 ( .INP(1'b1), .ZN(decodedPacket1_o[35]) );
  INVX0 U65 ( .INP(1'b1), .ZN(decodedPacket1_o[36]) );
  INVX0 U67 ( .INP(1'b1), .ZN(decodedPacket1_o[117]) );
  INVX0 U69 ( .INP(1'b1), .ZN(decodedPacket1_o[121]) );
  INVX0 U71 ( .INP(1'b1), .ZN(decodedPacket1_o[122]) );
  INVX0 U73 ( .INP(1'b1), .ZN(decodedPacket1_o[123]) );
  INVX0 U75 ( .INP(1'b1), .ZN(decodedPacket1_o[124]) );
  INVX0 U77 ( .INP(1'b1), .ZN(decodedPacket1_o[125]) );
  INVX0 U79 ( .INP(1'b1), .ZN(decodedPacket0_o[122]) );
  INVX0 U81 ( .INP(1'b1), .ZN(decodedPacket0_o[123]) );
  INVX0 U83 ( .INP(1'b1), .ZN(decodedPacket0_o[124]) );
  INVX0 U85 ( .INP(1'b1), .ZN(decodedPacket0_o[125]) );
  INVX0 U87 ( .INP(decodedPacket1_o[77]), .ZN(n316) );
  NBUFFX2 U88 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[73]) );
  NBUFFX2 U89 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[75]) );
  NBUFFX2 U90 ( .INP(decodedPacket1_o[76]), .Z(decodedPacket1_o[115]) );
  NBUFFX2 U91 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[69]) );
  NBUFFX2 U92 ( .INP(n511), .Z(decodedPacket1_o[76]) );
  NBUFFX2 U93 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[98]) );
  NBUFFX2 U94 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[118]) );
  NBUFFX2 U95 ( .INP(n511), .Z(decodedPacket1_o[74]) );
  NBUFFX2 U96 ( .INP(n511), .Z(decodedPacket1_o[77]) );
  NOR2X0 U97 ( .IN1(n506), .IN2(n459), .QN(n511) );
  INVX0 U98 ( .INP(n499), .ZN(n322) );
  NOR2X0 U99 ( .IN1(n336), .IN2(n308), .QN(decodedPacket1_o_119) );
  INVX0 U100 ( .INP(n482), .ZN(decodedPacket0_o[84]) );
  INVX0 U101 ( .INP(n509), .ZN(decodedPacket1_o[71]) );
  INVX0 U102 ( .INP(n468), .ZN(n317) );
  INVX0 U103 ( .INP(n500), .ZN(n318) );
  NOR2X0 U104 ( .IN1(n308), .IN2(n317), .QN(n472) );
  INVX0 U105 ( .INP(n460), .ZN(n321) );
  NAND2X1 U106 ( .IN1(n343), .IN2(n337), .QN(n489) );
  INVX0 U107 ( .INP(n423), .ZN(n334) );
  INVX0 U108 ( .INP(n485), .ZN(n323) );
  INVX0 U109 ( .INP(n412), .ZN(n338) );
  INVX0 U110 ( .INP(n467), .ZN(n319) );
  INVX0 U111 ( .INP(n463), .ZN(n320) );
  NOR2X0 U112 ( .IN1(n422), .IN2(n333), .QN(n455) );
  INVX0 U113 ( .INP(n424), .ZN(n333) );
  NAND2X1 U114 ( .IN1(n345), .IN2(n325), .QN(n456) );
  INVX0 U115 ( .INP(n478), .ZN(n326) );
  INVX0 U116 ( .INP(n443), .ZN(n325) );
  NOR2X0 U117 ( .IN1(n307), .IN2(n322), .QN(decodedPacket1_o[72]) );
  NOR2X0 U118 ( .IN1(n308), .IN2(n455), .QN(decodedPacket1_o_118) );
  NAND2X1 U119 ( .IN1(n315), .IN2(n395), .QN(n402) );
  NAND2X1 U120 ( .IN1(n315), .IN2(n481), .QN(n482) );
  INVX0 U121 ( .INP(n506), .ZN(n315) );
  NOR2X0 U122 ( .IN1(n412), .IN2(n405), .QN(n378) );
  NOR4X0 U123 ( .IN1(n464), .IN2(n463), .IN3(n478), .IN4(n462), .QN(n465) );
  NOR2X0 U124 ( .IN1(n307), .IN2(n424), .QN(decodedPacket1_o_120) );
  INVX0 U125 ( .INP(n399), .ZN(n337) );
  NOR2X0 U126 ( .IN1(n420), .IN2(n307), .QN(decodedPacket0_o[117]) );
  INVX0 U127 ( .INP(n417), .ZN(n332) );
  INVX0 U128 ( .INP(n442), .ZN(n343) );
  NOR2X0 U129 ( .IN1(n440), .IN2(n399), .QN(n412) );
  NOR2X0 U130 ( .IN1(n416), .IN2(n307), .QN(decodedPacket0_o[116]) );
  NOR4X0 U131 ( .IN1(n415), .IN2(n414), .IN3(n425), .IN4(n423), .QN(n416) );
  NOR2X0 U132 ( .IN1(n487), .IN2(n307), .QN(decodedPacket0_o[91]) );
  NOR4X0 U133 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(n487) );
  OR2X1 U134 ( .IN1(decodedPacket1_o[118]), .IN2(n224), .Q(
        decodedPacket0_o[118]) );
  AOI21X1 U135 ( .IN1(n335), .IN2(n421), .IN3(n308), .QN(n224) );
  INVX0 U136 ( .INP(n372), .ZN(n349) );
  INVX0 U137 ( .INP(n422), .ZN(n336) );
  NOR2X0 U138 ( .IN1(n474), .IN2(n308), .QN(n471) );
  NOR2X0 U139 ( .IN1(n343), .IN2(n346), .QN(n426) );
  OA21X1 U140 ( .IN1(n395), .IN2(n328), .IN3(n315), .Q(decodedPacket0_o[98])
         );
  INVX0 U141 ( .INP(n474), .ZN(n328) );
  NAND2X1 U142 ( .IN1(n406), .IN2(n335), .QN(n423) );
  INVX0 U143 ( .INP(n405), .ZN(n335) );
  INVX0 U144 ( .INP(n492), .ZN(n339) );
  NAND2X1 U145 ( .IN1(n315), .IN2(n457), .QN(n509) );
  NOR2X0 U146 ( .IN1(n350), .IN2(n345), .QN(n428) );
  INVX0 U147 ( .INP(n425), .ZN(n331) );
  NAND2X1 U148 ( .IN1(n473), .IN2(n474), .QN(n467) );
  INVX0 U149 ( .INP(n484), .ZN(n327) );
  INVX0 U150 ( .INP(n396), .ZN(n345) );
  NOR2X0 U151 ( .IN1(n403), .IN2(n376), .QN(n422) );
  INVX0 U152 ( .INP(n385), .ZN(n346) );
  NOR2X0 U153 ( .IN1(n443), .IN2(n403), .QN(n478) );
  NAND2X1 U154 ( .IN1(n346), .IN2(n377), .QN(n424) );
  NAND2X1 U155 ( .IN1(n380), .IN2(n342), .QN(n443) );
  NAND2X1 U156 ( .IN1(n375), .IN2(n354), .QN(n441) );
  INVX0 U157 ( .INP(n462), .ZN(n330) );
  NAND2X1 U158 ( .IN1(n349), .IN2(n377), .QN(n371) );
  NOR2X0 U159 ( .IN1(n441), .IN2(n376), .QN(n405) );
  NOR2X0 U274 ( .IN1(n442), .IN2(n376), .QN(n418) );
  NOR2X0 U298 ( .IN1(n396), .IN2(n376), .QN(n419) );
  NOR2X0 U333 ( .IN1(n400), .IN2(n399), .QN(n492) );
  NOR2X0 U334 ( .IN1(n370), .IN2(n402), .QN(decodedPacket0_o[107]) );
  NOR2X0 U335 ( .IN1(n369), .IN2(n402), .QN(decodedPacket0_o[108]) );
  NOR2X0 U336 ( .IN1(n368), .IN2(n402), .QN(decodedPacket0_o[109]) );
  NOR2X0 U337 ( .IN1(n367), .IN2(n402), .QN(decodedPacket0_o[110]) );
  NOR2X0 U338 ( .IN1(n366), .IN2(n402), .QN(decodedPacket0_o[111]) );
  NAND2X1 U339 ( .IN1(n476), .IN2(n386), .QN(n474) );
  NOR2X0 U340 ( .IN1(n362), .IN2(n482), .QN(decodedPacket0_o[85]) );
  NOR2X0 U341 ( .IN1(n361), .IN2(n482), .QN(decodedPacket0_o[86]) );
  NOR2X0 U342 ( .IN1(n360), .IN2(n482), .QN(decodedPacket0_o[87]) );
  NOR2X0 U343 ( .IN1(n359), .IN2(n482), .QN(decodedPacket0_o[88]) );
  NOR2X0 U344 ( .IN1(n358), .IN2(n482), .QN(decodedPacket0_o[89]) );
  NOR2X0 U345 ( .IN1(n357), .IN2(n482), .QN(decodedPacket0_o[90]) );
  NAND2X1 U346 ( .IN1(n316), .IN2(n342), .QN(decodedPacket0_o[73]) );
  NAND2X1 U347 ( .IN1(n316), .IN2(n341), .QN(decodedPacket0_o[74]) );
  NAND2X1 U348 ( .IN1(n316), .IN2(n340), .QN(decodedPacket0_o[75]) );
  NAND2X1 U349 ( .IN1(n316), .IN2(n329), .QN(decodedPacket0_o[76]) );
  NOR2X0 U350 ( .IN1(n475), .IN2(n308), .QN(decodedPacket0_o[83]) );
  NOR2X0 U351 ( .IN1(n496), .IN2(n307), .QN(decodedPacket0_o[94]) );
  NOR2X0 U352 ( .IN1(n497), .IN2(n308), .QN(decodedPacket0_o[95]) );
  NOR2X0 U353 ( .IN1(n494), .IN2(n308), .QN(decodedPacket0_o[92]) );
  NOR2X0 U354 ( .IN1(n492), .IN2(n503), .QN(n493) );
  NOR2X0 U355 ( .IN1(n498), .IN2(n307), .QN(decodedPacket0_o[96]) );
  NOR2X0 U356 ( .IN1(n470), .IN2(n308), .QN(decodedPacket0_o[78]) );
  NOR2X0 U357 ( .IN1(n495), .IN2(n308), .QN(decodedPacket0_o[93]) );
  INVX0 U358 ( .INP(n400), .ZN(n348) );
  NAND2X1 U359 ( .IN1(n509), .IN2(n352), .QN(decodedPacket0_o[71]) );
  NOR2X0 U360 ( .IN1(n316), .IN2(n356), .QN(decodedPacket1_o[78]) );
  NOR2X0 U361 ( .IN1(n316), .IN2(n355), .QN(decodedPacket1_o[83]) );
  NOR2X0 U362 ( .IN1(n436), .IN2(n427), .QN(n502) );
  INVX0 U363 ( .INP(n410), .ZN(n350) );
  NOR2X0 U364 ( .IN1(n352), .IN2(n443), .QN(n445) );
  NAND2X1 U365 ( .IN1(n444), .IN2(n352), .QN(n440) );
  NAND2X1 U366 ( .IN1(n348), .IN2(n377), .QN(n417) );
  NAND2X1 U367 ( .IN1(n343), .IN2(n377), .QN(n421) );
  NAND2X1 U368 ( .IN1(n476), .IN2(n344), .QN(n429) );
  NOR2X0 U369 ( .IN1(n503), .IN2(n502), .QN(n430) );
  INVX0 U370 ( .INP(n428), .ZN(n344) );
  NOR2X0 U371 ( .IN1(n501), .IN2(n357), .QN(n504) );
  NAND2X1 U372 ( .IN1(n350), .IN2(n476), .QN(n383) );
  NAND2X1 U373 ( .IN1(n476), .IN2(n345), .QN(n477) );
  INVX0 U374 ( .INP(n436), .ZN(n351) );
  NAND2X1 U375 ( .IN1(n337), .IN2(n411), .QN(n413) );
  INVX0 U376 ( .INP(n427), .ZN(n324) );
  NOR2X0 U377 ( .IN1(n352), .IN2(n450), .QN(n381) );
  NBUFFX2 U378 ( .INP(instPacketValid_i), .Z(decodedPacket0Valid_o) );
  NOR2X0 U379 ( .IN1(n352), .IN2(instPacket_i[104]), .QN(n379) );
  NAND2X1 U380 ( .IN1(n375), .IN2(instPacket_i[101]), .QN(n403) );
  INVX0 U381 ( .INP(instPacket_i[103]), .ZN(n352) );
  INVX0 U382 ( .INP(instPacket_i[101]), .ZN(n354) );
  INVX0 U383 ( .INP(instPacket_i[105]), .ZN(n342) );
  INVX0 U384 ( .INP(instPacket_i[102]), .ZN(n353) );
  INVX0 U385 ( .INP(instPacket_i[106]), .ZN(n341) );
  NOR2X0 U386 ( .IN1(instPacket_i[108]), .IN2(instPacket_i[107]), .QN(n374) );
  INVX0 U387 ( .INP(instPacket_i[108]), .ZN(n329) );
  NOR4X0 U388 ( .IN1(n390), .IN2(instPacket_i[127]), .IN3(instPacket_i[129]), 
        .IN4(instPacket_i[128]), .QN(n391) );
  NOR4X0 U389 ( .IN1(n389), .IN2(instPacket_i[121]), .IN3(instPacket_i[123]), 
        .IN4(instPacket_i[122]), .QN(n392) );
  NOR4X0 U390 ( .IN1(n387), .IN2(instPacket_i[109]), .IN3(instPacket_i[111]), 
        .IN4(instPacket_i[110]), .QN(n394) );
  NOR4X0 U391 ( .IN1(n388), .IN2(instPacket_i[115]), .IN3(instPacket_i[117]), 
        .IN4(instPacket_i[116]), .QN(n393) );
  NOR4X0 U392 ( .IN1(n483), .IN2(n484), .IN3(n307), .IN4(n452), .QN(n453) );
  NOR2X0 U393 ( .IN1(n365), .IN2(n402), .QN(decodedPacket0_o[112]) );
  INVX0 U394 ( .INP(instPacket_i_82), .ZN(n365) );
  NOR2X0 U395 ( .IN1(n364), .IN2(n402), .QN(decodedPacket0_o[113]) );
  INVX0 U396 ( .INP(instPacket_i_83), .ZN(n364) );
  NOR2X0 U397 ( .IN1(n363), .IN2(n402), .QN(decodedPacket0_o[114]) );
  INVX0 U398 ( .INP(instPacket_i_84), .ZN(n363) );
  INVX0 U399 ( .INP(n447), .ZN(n347) );
  NOR2X0 U400 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[102]), .QN(n448) );
  NOR2X0 U401 ( .IN1(n507), .IN2(n307), .QN(decodedPacket0_o[97]) );
  NOR4X0 U402 ( .IN1(n505), .IN2(n504), .IN3(n503), .IN4(n502), .QN(n507) );
  NOR2X0 U403 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[103]), .QN(n447) );
  INVX0 U404 ( .INP(instPacket_i_71), .ZN(N287) );
  XNOR2X1 U405 ( .IN1(n225), .IN2(instPacket_i_84), .Q(N300) );
  NAND2X1 U406 ( .IN1(instPacket_i_83), .IN2(\r340/carry[14] ), .QN(n225) );
  NBUFFX2 U407 ( .INP(instPacket_i[0]), .Z(decodedPacket0_o[0]) );
  NBUFFX2 U408 ( .INP(instPacket_i[1]), .Z(decodedPacket0_o[1]) );
  NBUFFX2 U409 ( .INP(instPacket_i[2]), .Z(decodedPacket0_o[2]) );
  NBUFFX2 U410 ( .INP(instPacket_i[3]), .Z(decodedPacket0_o[3]) );
  NBUFFX2 U411 ( .INP(instPacket_i[4]), .Z(decodedPacket0_o[4]) );
  NBUFFX2 U412 ( .INP(instPacket_i[37]), .Z(decodedPacket0_o[37]) );
  NBUFFX2 U413 ( .INP(instPacket_i[38]), .Z(decodedPacket0_o[38]) );
  NBUFFX2 U414 ( .INP(instPacket_i[39]), .Z(decodedPacket0_o[39]) );
  NBUFFX2 U415 ( .INP(instPacket_i[40]), .Z(decodedPacket0_o[40]) );
  NBUFFX2 U416 ( .INP(instPacket_i[41]), .Z(decodedPacket0_o[41]) );
  NBUFFX2 U417 ( .INP(instPacket_i[42]), .Z(decodedPacket0_o[42]) );
  NBUFFX2 U418 ( .INP(instPacket_i[43]), .Z(decodedPacket0_o[43]) );
  NBUFFX2 U419 ( .INP(instPacket_i[44]), .Z(decodedPacket0_o[44]) );
  NBUFFX2 U420 ( .INP(instPacket_i[45]), .Z(decodedPacket0_o[45]) );
  NBUFFX2 U421 ( .INP(instPacket_i[46]), .Z(decodedPacket0_o[46]) );
  NBUFFX2 U422 ( .INP(instPacket_i[47]), .Z(decodedPacket0_o[47]) );
  NBUFFX2 U423 ( .INP(instPacket_i[48]), .Z(decodedPacket0_o[48]) );
  NBUFFX2 U424 ( .INP(instPacket_i[49]), .Z(decodedPacket0_o[49]) );
  NBUFFX2 U425 ( .INP(instPacket_i[50]), .Z(decodedPacket0_o[50]) );
  NBUFFX2 U426 ( .INP(instPacket_i[51]), .Z(decodedPacket0_o[51]) );
  NBUFFX2 U427 ( .INP(instPacket_i[52]), .Z(decodedPacket0_o[52]) );
  NBUFFX2 U428 ( .INP(instPacket_i[53]), .Z(decodedPacket0_o[53]) );
  NBUFFX2 U429 ( .INP(instPacket_i[54]), .Z(decodedPacket0_o[54]) );
  NBUFFX2 U430 ( .INP(instPacket_i[55]), .Z(decodedPacket0_o[55]) );
  NBUFFX2 U431 ( .INP(instPacket_i[56]), .Z(decodedPacket0_o[56]) );
  NBUFFX2 U432 ( .INP(instPacket_i[57]), .Z(decodedPacket0_o[57]) );
  NBUFFX2 U433 ( .INP(instPacket_i[58]), .Z(decodedPacket0_o[58]) );
  NBUFFX2 U434 ( .INP(instPacket_i[59]), .Z(decodedPacket0_o[59]) );
  NBUFFX2 U435 ( .INP(instPacket_i[60]), .Z(decodedPacket0_o[60]) );
  NBUFFX2 U436 ( .INP(instPacket_i[61]), .Z(decodedPacket0_o[61]) );
  NBUFFX2 U437 ( .INP(instPacket_i[62]), .Z(decodedPacket0_o[62]) );
  NBUFFX2 U438 ( .INP(instPacket_i[63]), .Z(decodedPacket0_o[63]) );
  NBUFFX2 U439 ( .INP(instPacket_i[64]), .Z(decodedPacket0_o[64]) );
  NBUFFX2 U440 ( .INP(instPacket_i[65]), .Z(decodedPacket0_o[65]) );
  NBUFFX2 U441 ( .INP(instPacket_i[66]), .Z(decodedPacket0_o[66]) );
  NBUFFX2 U442 ( .INP(instPacket_i[67]), .Z(decodedPacket0_o[67]) );
  NBUFFX2 U443 ( .INP(instPacket_i[68]), .Z(decodedPacket0_o[68]) );
  NAND2X1 U444 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[104]), .QN(n450)
         );
  NBUFFX2 U445 ( .INP(instPacket_i[0]), .Z(decodedPacket1_o[0]) );
  NBUFFX2 U446 ( .INP(instPacket_i[1]), .Z(decodedPacket1_o[1]) );
  NBUFFX2 U447 ( .INP(instPacket_i[2]), .Z(decodedPacket1_o[2]) );
  NBUFFX2 U448 ( .INP(instPacket_i[3]), .Z(decodedPacket1_o[3]) );
  NBUFFX2 U449 ( .INP(instPacket_i[4]), .Z(decodedPacket1_o[4]) );
  NBUFFX2 U450 ( .INP(instPacket_i[37]), .Z(decodedPacket1_o[37]) );
  NBUFFX2 U451 ( .INP(instPacket_i[38]), .Z(decodedPacket1_o[38]) );
  NBUFFX2 U452 ( .INP(instPacket_i[39]), .Z(decodedPacket1_o[39]) );
  NBUFFX2 U453 ( .INP(instPacket_i[40]), .Z(decodedPacket1_o[40]) );
  NBUFFX2 U454 ( .INP(instPacket_i[41]), .Z(decodedPacket1_o[41]) );
  NBUFFX2 U455 ( .INP(instPacket_i[42]), .Z(decodedPacket1_o[42]) );
  NBUFFX2 U456 ( .INP(instPacket_i[43]), .Z(decodedPacket1_o[43]) );
  NBUFFX2 U457 ( .INP(instPacket_i[44]), .Z(decodedPacket1_o[44]) );
  NBUFFX2 U458 ( .INP(instPacket_i[45]), .Z(decodedPacket1_o[45]) );
  NBUFFX2 U459 ( .INP(instPacket_i[46]), .Z(decodedPacket1_o[46]) );
  NBUFFX2 U460 ( .INP(instPacket_i[47]), .Z(decodedPacket1_o[47]) );
  NBUFFX2 U461 ( .INP(instPacket_i[48]), .Z(decodedPacket1_o[48]) );
  NBUFFX2 U462 ( .INP(instPacket_i[49]), .Z(decodedPacket1_o[49]) );
  NBUFFX2 U463 ( .INP(instPacket_i[50]), .Z(decodedPacket1_o[50]) );
  NBUFFX2 U464 ( .INP(instPacket_i[51]), .Z(decodedPacket1_o[51]) );
  NBUFFX2 U465 ( .INP(instPacket_i[52]), .Z(decodedPacket1_o[52]) );
  NBUFFX2 U466 ( .INP(instPacket_i[53]), .Z(decodedPacket1_o[53]) );
  NBUFFX2 U467 ( .INP(instPacket_i[54]), .Z(decodedPacket1_o[54]) );
  NBUFFX2 U468 ( .INP(instPacket_i[55]), .Z(decodedPacket1_o[55]) );
  NBUFFX2 U469 ( .INP(instPacket_i[56]), .Z(decodedPacket1_o[56]) );
  NBUFFX2 U470 ( .INP(instPacket_i[57]), .Z(decodedPacket1_o[57]) );
  NBUFFX2 U471 ( .INP(instPacket_i[58]), .Z(decodedPacket1_o[58]) );
  NBUFFX2 U472 ( .INP(instPacket_i[59]), .Z(decodedPacket1_o[59]) );
  NBUFFX2 U473 ( .INP(instPacket_i[60]), .Z(decodedPacket1_o[60]) );
  NBUFFX2 U474 ( .INP(instPacket_i[61]), .Z(decodedPacket1_o[61]) );
  NBUFFX2 U475 ( .INP(instPacket_i[62]), .Z(decodedPacket1_o[62]) );
  NBUFFX2 U476 ( .INP(instPacket_i[63]), .Z(decodedPacket1_o[63]) );
  NBUFFX2 U477 ( .INP(instPacket_i[64]), .Z(decodedPacket1_o[64]) );
  NBUFFX2 U478 ( .INP(instPacket_i[65]), .Z(decodedPacket1_o[65]) );
  NBUFFX2 U479 ( .INP(instPacket_i[66]), .Z(decodedPacket1_o[66]) );
  NBUFFX2 U480 ( .INP(instPacket_i[67]), .Z(decodedPacket1_o[67]) );
  NBUFFX2 U481 ( .INP(instPacket_i[68]), .Z(decodedPacket1_o[68]) );
  NOR2X0 U482 ( .IN1(n450), .IN2(instPacket_i[101]), .QN(n444) );
  INVX0 U483 ( .INP(instPacket_i[107]), .ZN(n340) );
  INVX0 U484 ( .INP(instPacket_i_90), .ZN(n357) );
  NAND2X1 U485 ( .IN1(n325), .IN2(instPacket_i[101]), .QN(n427) );
  NOR2X0 U486 ( .IN1(n437), .IN2(n354), .QN(n438) );
  INVX0 U487 ( .INP(instPacket_i_85), .ZN(n362) );
  INVX0 U488 ( .INP(instPacket_i_93), .ZN(n356) );
  INVX0 U489 ( .INP(instPacket_i_98), .ZN(n355) );
  INVX0 U490 ( .INP(instPacket_i_77), .ZN(n370) );
  INVX0 U491 ( .INP(instPacket_i_78), .ZN(n369) );
  INVX0 U492 ( .INP(instPacket_i_79), .ZN(n368) );
  INVX0 U493 ( .INP(instPacket_i_80), .ZN(n367) );
  INVX0 U494 ( .INP(instPacket_i_81), .ZN(n366) );
  INVX0 U495 ( .INP(instPacket_i_86), .ZN(n361) );
  INVX0 U496 ( .INP(instPacket_i_87), .ZN(n360) );
  INVX0 U497 ( .INP(instPacket_i_88), .ZN(n359) );
  INVX0 U498 ( .INP(instPacket_i_89), .ZN(n358) );
  NBUFFX2 U499 ( .INP(n508), .Z(n312) );
  NBUFFX2 U500 ( .INP(n510), .Z(decodedPacket0_o[121]) );
  NBUFFX2 U501 ( .INP(n510), .Z(n314) );
  NAND4X0 U502 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n307) );
  NAND4X0 U503 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n308) );
  XOR2X1 U504 ( .IN1(\r340/carry[14] ), .IN2(instPacket_i_83), .Q(N299) );
  AND2X1 U505 ( .IN1(instPacket_i_82), .IN2(\r340/carry[13] ), .Q(
        \r340/carry[14] ) );
  XOR2X1 U506 ( .IN1(\r340/carry[13] ), .IN2(instPacket_i_82), .Q(N298) );
  AND2X1 U507 ( .IN1(instPacket_i_81), .IN2(\r340/carry[12] ), .Q(
        \r340/carry[13] ) );
  XOR2X1 U508 ( .IN1(\r340/carry[12] ), .IN2(instPacket_i_81), .Q(N297) );
  AND2X1 U509 ( .IN1(instPacket_i_80), .IN2(\r340/carry[11] ), .Q(
        \r340/carry[12] ) );
  XOR2X1 U510 ( .IN1(\r340/carry[11] ), .IN2(instPacket_i_80), .Q(N296) );
  AND2X1 U511 ( .IN1(instPacket_i_79), .IN2(\r340/carry[10] ), .Q(
        \r340/carry[11] ) );
  XOR2X1 U512 ( .IN1(\r340/carry[10] ), .IN2(instPacket_i_79), .Q(N295) );
  AND2X1 U513 ( .IN1(instPacket_i_78), .IN2(\r340/carry[9] ), .Q(
        \r340/carry[10] ) );
  XOR2X1 U514 ( .IN1(\r340/carry[9] ), .IN2(instPacket_i_78), .Q(N294) );
  AND2X1 U515 ( .IN1(instPacket_i_77), .IN2(\r340/carry[8] ), .Q(
        \r340/carry[9] ) );
  XOR2X1 U516 ( .IN1(\r340/carry[8] ), .IN2(instPacket_i_77), .Q(N293) );
  AND2X1 U517 ( .IN1(instPacket_i_76), .IN2(\r340/carry[7] ), .Q(
        \r340/carry[8] ) );
  XOR2X1 U518 ( .IN1(\r340/carry[7] ), .IN2(instPacket_i_76), .Q(N292) );
  AND2X1 U519 ( .IN1(instPacket_i_75), .IN2(\r340/carry[6] ), .Q(
        \r340/carry[7] ) );
  XOR2X1 U520 ( .IN1(\r340/carry[6] ), .IN2(instPacket_i_75), .Q(N291) );
  AND2X1 U521 ( .IN1(instPacket_i_74), .IN2(\r340/carry[5] ), .Q(
        \r340/carry[6] ) );
  XOR2X1 U522 ( .IN1(\r340/carry[5] ), .IN2(instPacket_i_74), .Q(N290) );
  AND2X1 U523 ( .IN1(instPacket_i_73), .IN2(\r340/carry[4] ), .Q(
        \r340/carry[5] ) );
  XOR2X1 U524 ( .IN1(\r340/carry[4] ), .IN2(instPacket_i_73), .Q(N289) );
  AND2X1 U525 ( .IN1(instPacket_i_72), .IN2(instPacket_i_71), .Q(
        \r340/carry[4] ) );
  XOR2X1 U526 ( .IN1(instPacket_i_71), .IN2(instPacket_i_72), .Q(N288) );
  XOR2X1 U527 ( .IN1(\r339/carry[5] ), .IN2(instPacket_i_90), .Q(N284) );
endmodule


module Decode_PISA_1 ( instPacketValid_i, instPacket_i, decodedPacket0Valid_o, 
        decodedPacket0_o, decodedPacket1Valid_o, decodedPacket1_o );
  input [132:0] instPacket_i;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  input instPacketValid_i;
  output decodedPacket0Valid_o, decodedPacket1Valid_o;
  wire   instPacket_i_98, instPacket_i_97, instPacket_i_96, instPacket_i_95,
         instPacket_i_94, instPacket_i_93, instPacket_i_92, instPacket_i_91,
         instPacket_i_90, instPacket_i_89, instPacket_i_88, instPacket_i_87,
         instPacket_i_86, instPacket_i_85, instPacket_i_84, instPacket_i_83,
         instPacket_i_82, instPacket_i_81, instPacket_i_80, instPacket_i_79,
         instPacket_i_78, instPacket_i_77, instPacket_i_76, instPacket_i_75,
         instPacket_i_74, instPacket_i_73, instPacket_i_72, instPacket_i_71,
         instPacket_i_36, instPacket_i_35, instPacket_i_34, instPacket_i_33,
         instPacket_i_32, instPacket_i_31, instPacket_i_30, instPacket_i_29,
         instPacket_i_28, instPacket_i_27, instPacket_i_26, instPacket_i_25,
         instPacket_i_24, instPacket_i_23, instPacket_i_22, instPacket_i_21,
         instPacket_i_20, instPacket_i_19, instPacket_i_18, instPacket_i_17,
         instPacket_i_16, instPacket_i_15, instPacket_i_14, instPacket_i_13,
         instPacket_i_12, instPacket_i_11, instPacket_i_10, instPacket_i_9,
         instPacket_i_8, instPacket_i_7, instPacket_i_6, instPacket_i_5, n510,
         decodedPacket1_o_120, decodedPacket1_o_119, decodedPacket1_o_118,
         n511, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         \r340/carry[14] , \r340/carry[13] , \r340/carry[12] ,
         \r340/carry[11] , \r340/carry[10] , \r340/carry[9] , \r340/carry[8] ,
         \r340/carry[7] , \r340/carry[6] , \r340/carry[5] , \r340/carry[4] ,
         \r339/carry[5] , \r339/carry[4] , \r339/carry[3] , \r339/carry[2] ,
         n224, n225, n307, n308, n312, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509;
  assign instPacket_i_98 = instPacket_i[98];
  assign instPacket_i_97 = instPacket_i[97];
  assign instPacket_i_96 = instPacket_i[96];
  assign instPacket_i_95 = instPacket_i[95];
  assign instPacket_i_94 = instPacket_i[94];
  assign instPacket_i_93 = instPacket_i[93];
  assign instPacket_i_92 = instPacket_i[92];
  assign instPacket_i_91 = instPacket_i[91];
  assign instPacket_i_90 = instPacket_i[90];
  assign instPacket_i_89 = instPacket_i[89];
  assign instPacket_i_88 = instPacket_i[88];
  assign instPacket_i_87 = instPacket_i[87];
  assign instPacket_i_86 = instPacket_i[86];
  assign instPacket_i_85 = instPacket_i[85];
  assign instPacket_i_84 = instPacket_i[84];
  assign instPacket_i_83 = instPacket_i[83];
  assign instPacket_i_82 = instPacket_i[82];
  assign instPacket_i_81 = instPacket_i[81];
  assign instPacket_i_80 = instPacket_i[80];
  assign instPacket_i_79 = instPacket_i[79];
  assign instPacket_i_78 = instPacket_i[78];
  assign instPacket_i_77 = instPacket_i[77];
  assign instPacket_i_76 = instPacket_i[76];
  assign instPacket_i_75 = instPacket_i[75];
  assign instPacket_i_74 = instPacket_i[74];
  assign instPacket_i_73 = instPacket_i[73];
  assign instPacket_i_72 = instPacket_i[72];
  assign instPacket_i_71 = instPacket_i[71];
  assign instPacket_i_36 = instPacket_i[36];
  assign instPacket_i_35 = instPacket_i[35];
  assign instPacket_i_34 = instPacket_i[34];
  assign instPacket_i_33 = instPacket_i[33];
  assign instPacket_i_32 = instPacket_i[32];
  assign instPacket_i_31 = instPacket_i[31];
  assign instPacket_i_30 = instPacket_i[30];
  assign instPacket_i_29 = instPacket_i[29];
  assign instPacket_i_28 = instPacket_i[28];
  assign instPacket_i_27 = instPacket_i[27];
  assign instPacket_i_26 = instPacket_i[26];
  assign instPacket_i_25 = instPacket_i[25];
  assign instPacket_i_24 = instPacket_i[24];
  assign instPacket_i_23 = instPacket_i[23];
  assign instPacket_i_22 = instPacket_i[22];
  assign instPacket_i_21 = instPacket_i[21];
  assign instPacket_i_20 = instPacket_i[20];
  assign instPacket_i_19 = instPacket_i[19];
  assign instPacket_i_18 = instPacket_i[18];
  assign instPacket_i_17 = instPacket_i[17];
  assign instPacket_i_16 = instPacket_i[16];
  assign instPacket_i_15 = instPacket_i[15];
  assign instPacket_i_14 = instPacket_i[14];
  assign instPacket_i_13 = instPacket_i[13];
  assign instPacket_i_12 = instPacket_i[12];
  assign instPacket_i_11 = instPacket_i[11];
  assign instPacket_i_10 = instPacket_i[10];
  assign instPacket_i_9 = instPacket_i[9];
  assign instPacket_i_8 = instPacket_i[8];
  assign instPacket_i_7 = instPacket_i[7];
  assign instPacket_i_6 = instPacket_i[6];
  assign instPacket_i_5 = instPacket_i[5];
  assign decodedPacket1_o[120] = decodedPacket1_o_120;
  assign decodedPacket1_o[119] = decodedPacket1_o_119;
  assign decodedPacket1_o[116] = decodedPacket1_o_118;
  assign N285 = instPacket_i[69];
  assign N286 = instPacket_i[70];

  AND2X1 U160 ( .IN1(N285), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[99]) );
  AO21X1 U161 ( .IN1(N284), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[97]) );
  AND2X1 U162 ( .IN1(decodedPacket1_o_119), .IN2(N283), .Q(
        decodedPacket1_o[96]) );
  AND2X1 U163 ( .IN1(decodedPacket1_o_119), .IN2(N282), .Q(
        decodedPacket1_o[95]) );
  AND2X1 U164 ( .IN1(decodedPacket1_o_119), .IN2(N281), .Q(
        decodedPacket1_o[94]) );
  AND2X1 U165 ( .IN1(decodedPacket1_o_119), .IN2(N280), .Q(
        decodedPacket1_o[93]) );
  AO21X1 U166 ( .IN1(n362), .IN2(decodedPacket1_o_119), .IN3(
        decodedPacket1_o[72]), .Q(decodedPacket1_o[92]) );
  OR2X1 U167 ( .IN1(decodedPacket1_o_119), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[91]) );
  AO22X1 U168 ( .IN1(decodedPacket1_o_120), .IN2(N284), .IN3(instPacket_i_90), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[90]) );
  AO22X1 U169 ( .IN1(decodedPacket1_o_120), .IN2(N283), .IN3(instPacket_i_89), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[89]) );
  AO22X1 U170 ( .IN1(decodedPacket1_o_120), .IN2(N282), .IN3(instPacket_i_88), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[88]) );
  AO22X1 U171 ( .IN1(decodedPacket1_o_120), .IN2(N281), .IN3(instPacket_i_87), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[87]) );
  AO22X1 U172 ( .IN1(decodedPacket1_o_120), .IN2(N280), .IN3(instPacket_i_86), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[86]) );
  AO22X1 U173 ( .IN1(decodedPacket1_o_120), .IN2(n362), .IN3(instPacket_i_85), 
        .IN4(decodedPacket1_o[72]), .Q(decodedPacket1_o[85]) );
  OR2X1 U174 ( .IN1(decodedPacket1_o_120), .IN2(decodedPacket1_o[72]), .Q(
        decodedPacket1_o[84]) );
  AND2X1 U175 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_97), .Q(
        decodedPacket1_o[82]) );
  AND2X1 U176 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_96), .Q(
        decodedPacket1_o[81]) );
  AND2X1 U177 ( .IN1(decodedPacket1_o[77]), .IN2(instPacket_i_95), .Q(
        decodedPacket1_o[80]) );
  AND2X1 U178 ( .IN1(decodedPacket1_o[76]), .IN2(instPacket_i_94), .Q(
        decodedPacket1_o[79]) );
  AND2X1 U179 ( .IN1(N300), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[114]) );
  AND2X1 U180 ( .IN1(N299), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[113]) );
  AND2X1 U181 ( .IN1(N298), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[112]) );
  AND2X1 U182 ( .IN1(N297), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[111]) );
  AND2X1 U183 ( .IN1(N296), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[110]) );
  AND2X1 U184 ( .IN1(N295), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[109]) );
  AND2X1 U185 ( .IN1(N294), .IN2(decodedPacket1_o_118), .Q(
        decodedPacket1_o[108]) );
  AND2X1 U186 ( .IN1(N293), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[107]) );
  AND2X1 U187 ( .IN1(N292), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[106]) );
  AND2X1 U188 ( .IN1(N291), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[105]) );
  AND2X1 U189 ( .IN1(N290), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[104]) );
  AND2X1 U190 ( .IN1(N289), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[103]) );
  AND2X1 U191 ( .IN1(N288), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[102]) );
  AND2X1 U192 ( .IN1(N287), .IN2(decodedPacket1_o[118]), .Q(
        decodedPacket1_o[101]) );
  AND2X1 U193 ( .IN1(N286), .IN2(decodedPacket1_o[98]), .Q(
        decodedPacket1_o[100]) );
  AND2X1 U194 ( .IN1(instPacketValid_i), .IN2(decodedPacket1_o[76]), .Q(
        decodedPacket1Valid_o) );
  AO22X1 U195 ( .IN1(instPacket_i_9), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_73), .IN4(n312), .Q(decodedPacket0_o[9]) );
  AND2X1 U196 ( .IN1(decodedPacket0_o[98]), .IN2(N285), .Q(
        decodedPacket0_o[99]) );
  AO21X1 U197 ( .IN1(instPacket_i_82), .IN2(n500), .IN3(n499), .Q(n505) );
  OA221X1 U198 ( .IN1(n318), .IN2(n366), .IN3(n501), .IN4(n358), .IN5(n339), 
        .Q(n498) );
  OA221X1 U199 ( .IN1(n318), .IN2(n367), .IN3(n501), .IN4(n359), .IN5(n339), 
        .Q(n497) );
  OA221X1 U200 ( .IN1(n318), .IN2(n368), .IN3(n501), .IN4(n360), .IN5(n339), 
        .Q(n496) );
  OA221X1 U201 ( .IN1(n318), .IN2(n369), .IN3(n501), .IN4(n361), .IN5(n339), 
        .Q(n495) );
  OA221X1 U202 ( .IN1(n318), .IN2(n370), .IN3(n501), .IN4(n362), .IN5(n493), 
        .Q(n494) );
  AND3X1 U203 ( .IN1(n491), .IN2(n336), .IN3(n334), .Q(n501) );
  NAND4X0 U204 ( .IN1(n490), .IN2(n319), .IN3(n489), .IN4(n488), .QN(n500) );
  NAND4X0 U205 ( .IN1(n489), .IN2(n339), .IN3(n326), .IN4(n336), .QN(n486) );
  AO22X1 U206 ( .IN1(instPacket_i_8), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_72), .IN4(n508), .Q(decodedPacket0_o[8]) );
  NAND4X0 U207 ( .IN1(n490), .IN2(n331), .IN3(n323), .IN4(n480), .QN(n481) );
  NOR3X0 U208 ( .IN1(n479), .IN2(n333), .IN3(n478), .QN(n480) );
  OA21X1 U209 ( .IN1(n345), .IN2(n346), .IN3(n337), .Q(n479) );
  AND3X1 U210 ( .IN1(n477), .IN2(n320), .IN3(n327), .Q(n490) );
  OA221X1 U211 ( .IN1(n317), .IN2(n355), .IN3(n357), .IN4(n474), .IN5(n473), 
        .Q(n475) );
  AO22X1 U212 ( .IN1(n472), .IN2(instPacket_i_97), .IN3(n471), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[82]) );
  AO22X1 U213 ( .IN1(n472), .IN2(instPacket_i_96), .IN3(n471), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[81]) );
  AO22X1 U214 ( .IN1(n472), .IN2(instPacket_i_95), .IN3(n471), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[80]) );
  AO22X1 U215 ( .IN1(instPacket_i_7), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_71), .IN4(n508), .Q(decodedPacket0_o[7]) );
  AO22X1 U216 ( .IN1(n472), .IN2(instPacket_i_94), .IN3(n471), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[79]) );
  OA221X1 U217 ( .IN1(n317), .IN2(n356), .IN3(n362), .IN4(n474), .IN5(n469), 
        .Q(n470) );
  OA21X1 U218 ( .IN1(n467), .IN2(n468), .IN3(n315), .Q(decodedPacket0_o[77])
         );
  NAND4X0 U219 ( .IN1(n466), .IN2(n327), .IN3(n323), .IN4(n465), .QN(n468) );
  NAND3X0 U220 ( .IN1(n461), .IN2(n488), .IN3(n460), .QN(n485) );
  AO21X1 U221 ( .IN1(instPacket_i[104]), .IN2(n458), .IN3(decodedPacket1_o[72]), .Q(decodedPacket0_o[72]) );
  NAND3X0 U222 ( .IN1(n456), .IN2(n461), .IN3(n455), .QN(n457) );
  AO21X1 U223 ( .IN1(instPacket_i[102]), .IN2(n458), .IN3(decodedPacket1_o[70]), .Q(decodedPacket0_o[70]) );
  AO21X1 U224 ( .IN1(n315), .IN2(n321), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket1_o[70]) );
  AO22X1 U225 ( .IN1(instPacket_i_6), .IN2(decodedPacket0_o[121]), .IN3(N286), 
        .IN4(n508), .Q(decodedPacket0_o[6]) );
  AND2X1 U226 ( .IN1(n458), .IN2(instPacket_i[101]), .Q(decodedPacket0_o[69])
         );
  NAND4X0 U227 ( .IN1(n488), .IN2(n329), .IN3(n454), .IN4(n453), .QN(n458) );
  AND2X1 U228 ( .IN1(instPacket_i[106]), .IN2(n451), .Q(n452) );
  NAND4X0 U229 ( .IN1(n347), .IN2(n340), .IN3(n450), .IN4(n449), .QN(n451) );
  OA22X1 U230 ( .IN1(instPacket_i[105]), .IN2(n352), .IN3(n448), .IN4(n342), 
        .Q(n449) );
  AO22X1 U231 ( .IN1(n476), .IN2(n446), .IN3(n445), .IN4(n444), .Q(n484) );
  NAND4X0 U232 ( .IN1(n442), .IN2(n441), .IN3(n440), .IN4(n439), .QN(n446) );
  NOR3X0 U233 ( .IN1(n438), .IN2(n348), .IN3(n349), .QN(n439) );
  OA21X1 U234 ( .IN1(instPacket_i[103]), .IN2(n450), .IN3(n436), .Q(n437) );
  NAND4X0 U235 ( .IN1(n466), .IN2(n319), .IN3(n435), .IN4(n334), .QN(n483) );
  AND2X1 U236 ( .IN1(n320), .IN2(n434), .Q(n435) );
  OA21X1 U237 ( .IN1(n348), .IN2(n349), .IN3(n325), .Q(n463) );
  AND2X1 U238 ( .IN1(n469), .IN2(n433), .Q(n473) );
  NAND3X0 U239 ( .IN1(n325), .IN2(n354), .IN3(n351), .QN(n433) );
  OR2X1 U240 ( .IN1(n440), .IN2(n443), .Q(n469) );
  AND4X1 U241 ( .IN1(n432), .IN2(n431), .IN3(n430), .IN4(n429), .Q(n466) );
  NOR3X0 U242 ( .IN1(n450), .IN2(instPacket_i[103]), .IN3(n427), .QN(n503) );
  AOI22X1 U243 ( .IN1(n340), .IN2(n341), .IN3(instPacket_i[103]), .IN4(
        instPacket_i[104]), .QN(n454) );
  OR2X1 U244 ( .IN1(n443), .IN2(n426), .Q(n488) );
  AO22X1 U245 ( .IN1(instPacket_i_5), .IN2(decodedPacket0_o[121]), .IN3(N285), 
        .IN4(n508), .Q(decodedPacket0_o[5]) );
  AND2X1 U246 ( .IN1(instPacket_i_36), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[36]) );
  AND2X1 U247 ( .IN1(instPacket_i_35), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[35]) );
  AND2X1 U248 ( .IN1(instPacket_i_34), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[34]) );
  AND2X1 U249 ( .IN1(instPacket_i_33), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[33]) );
  AND2X1 U250 ( .IN1(instPacket_i_32), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[32]) );
  AND2X1 U251 ( .IN1(instPacket_i_31), .IN2(decodedPacket0_o[121]), .Q(
        decodedPacket0_o[31]) );
  AO22X1 U252 ( .IN1(instPacket_i_30), .IN2(decodedPacket0_o[121]), .IN3(n508), 
        .IN4(instPacket_i_94), .Q(decodedPacket0_o[30]) );
  AO22X1 U253 ( .IN1(instPacket_i_29), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_93), .Q(decodedPacket0_o[29]) );
  AO22X1 U254 ( .IN1(instPacket_i_28), .IN2(n314), .IN3(instPacket_i_92), 
        .IN4(n508), .Q(decodedPacket0_o[28]) );
  AO22X1 U255 ( .IN1(instPacket_i_27), .IN2(n510), .IN3(instPacket_i_91), 
        .IN4(n508), .Q(decodedPacket0_o[27]) );
  AO22X1 U256 ( .IN1(instPacket_i_26), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_90), .Q(decodedPacket0_o[26]) );
  AO22X1 U257 ( .IN1(instPacket_i_25), .IN2(n314), .IN3(n312), .IN4(
        instPacket_i_89), .Q(decodedPacket0_o[25]) );
  AO22X1 U258 ( .IN1(instPacket_i_24), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_88), .Q(decodedPacket0_o[24]) );
  AO22X1 U259 ( .IN1(instPacket_i_23), .IN2(n314), .IN3(n312), .IN4(
        instPacket_i_87), .Q(decodedPacket0_o[23]) );
  AO22X1 U260 ( .IN1(instPacket_i_22), .IN2(n510), .IN3(n508), .IN4(
        instPacket_i_86), .Q(decodedPacket0_o[22]) );
  AO22X1 U261 ( .IN1(instPacket_i_21), .IN2(n314), .IN3(n508), .IN4(
        instPacket_i_85), .Q(decodedPacket0_o[21]) );
  AO22X1 U262 ( .IN1(instPacket_i_20), .IN2(n510), .IN3(instPacket_i_84), 
        .IN4(n312), .Q(decodedPacket0_o[20]) );
  AO22X1 U263 ( .IN1(instPacket_i_19), .IN2(n314), .IN3(instPacket_i_83), 
        .IN4(n312), .Q(decodedPacket0_o[19]) );
  AO22X1 U264 ( .IN1(instPacket_i_18), .IN2(n510), .IN3(instPacket_i_82), 
        .IN4(n312), .Q(decodedPacket0_o[18]) );
  AO22X1 U265 ( .IN1(instPacket_i_17), .IN2(n314), .IN3(instPacket_i_81), 
        .IN4(n312), .Q(decodedPacket0_o[17]) );
  AO22X1 U266 ( .IN1(instPacket_i_16), .IN2(n314), .IN3(instPacket_i_80), 
        .IN4(n312), .Q(decodedPacket0_o[16]) );
  AO22X1 U267 ( .IN1(instPacket_i_15), .IN2(n314), .IN3(instPacket_i_79), 
        .IN4(n312), .Q(decodedPacket0_o[15]) );
  AO22X1 U268 ( .IN1(instPacket_i_14), .IN2(n314), .IN3(instPacket_i_78), 
        .IN4(n312), .Q(decodedPacket0_o[14]) );
  AO22X1 U269 ( .IN1(instPacket_i_13), .IN2(n314), .IN3(instPacket_i_77), 
        .IN4(n312), .Q(decodedPacket0_o[13]) );
  AO22X1 U270 ( .IN1(instPacket_i_12), .IN2(n314), .IN3(instPacket_i_76), 
        .IN4(n312), .Q(decodedPacket0_o[12]) );
  AO21X1 U271 ( .IN1(n315), .IN2(n425), .IN3(decodedPacket1_o_120), .Q(
        decodedPacket0_o[120]) );
  AO22X1 U272 ( .IN1(instPacket_i_11), .IN2(decodedPacket0_o[121]), .IN3(
        instPacket_i_75), .IN4(n312), .Q(decodedPacket0_o[11]) );
  AO21X1 U273 ( .IN1(n315), .IN2(n423), .IN3(decodedPacket1_o_119), .Q(
        decodedPacket0_o[119]) );
  NOR3X0 U275 ( .IN1(n419), .IN2(n332), .IN3(n418), .QN(n420) );
  NAND3X0 U276 ( .IN1(n413), .IN2(n338), .IN3(n455), .QN(n415) );
  NAND3X0 U277 ( .IN1(n426), .IN2(n410), .IN3(n409), .QN(n411) );
  AND2X1 U278 ( .IN1(n315), .IN2(n408), .Q(decodedPacket0_o[115]) );
  NAND4X0 U279 ( .IN1(n459), .IN2(n334), .IN3(n331), .IN4(n407), .QN(n408) );
  NAND4X0 U280 ( .IN1(n349), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n407) );
  AND2X1 U281 ( .IN1(n455), .IN2(n322), .Q(n459) );
  NAND3X0 U282 ( .IN1(n326), .IN2(n461), .IN3(n460), .QN(n499) );
  OA21X1 U283 ( .IN1(n441), .IN2(n443), .IN3(n456), .Q(n460) );
  OR2X1 U284 ( .IN1(n443), .IN2(n404), .Q(n461) );
  AO22X1 U285 ( .IN1(instPacket_i_10), .IN2(n314), .IN3(instPacket_i_74), 
        .IN4(n312), .Q(decodedPacket0_o[10]) );
  AND2X1 U286 ( .IN1(n315), .IN2(n414), .Q(n508) );
  AO21X1 U287 ( .IN1(n337), .IN2(n401), .IN3(n492), .Q(n414) );
  OA21X1 U288 ( .IN1(n464), .IN2(n412), .IN3(n315), .Q(n510) );
  AND2X1 U289 ( .IN1(n337), .IN2(n398), .Q(n464) );
  NAND4X0 U290 ( .IN1(n426), .IN2(n428), .IN3(n397), .IN4(n404), .QN(n398) );
  AND2X1 U291 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_76), .Q(
        decodedPacket0_o[106]) );
  AND2X1 U292 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_75), .Q(
        decodedPacket0_o[105]) );
  AND2X1 U293 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_74), .Q(
        decodedPacket0_o[104]) );
  AND2X1 U294 ( .IN1(instPacket_i_73), .IN2(decodedPacket0_o[98]), .Q(
        decodedPacket0_o[103]) );
  AND2X1 U295 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_72), .Q(
        decodedPacket0_o[102]) );
  AND2X1 U296 ( .IN1(decodedPacket0_o[98]), .IN2(instPacket_i_71), .Q(
        decodedPacket0_o[101]) );
  AND2X1 U297 ( .IN1(decodedPacket0_o[98]), .IN2(N286), .Q(
        decodedPacket0_o[100]) );
  NAND4X0 U299 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n506) );
  OR3X1 U300 ( .IN1(instPacket_i[132]), .IN2(instPacket_i[131]), .IN3(
        instPacket_i[130]), .Q(n390) );
  OR3X1 U301 ( .IN1(instPacket_i[126]), .IN2(instPacket_i[125]), .IN3(
        instPacket_i[124]), .Q(n389) );
  OR3X1 U302 ( .IN1(instPacket_i[120]), .IN2(instPacket_i[119]), .IN3(
        instPacket_i[118]), .Q(n388) );
  OR3X1 U303 ( .IN1(instPacket_i[114]), .IN2(instPacket_i[113]), .IN3(
        instPacket_i[112]), .Q(n387) );
  NAND3X0 U304 ( .IN1(n403), .IN2(n385), .IN3(n404), .QN(n386) );
  NAND3X0 U305 ( .IN1(n330), .IN2(n384), .IN3(n491), .QN(n395) );
  AND4X1 U306 ( .IN1(n432), .IN2(n431), .IN3(n383), .IN4(n434), .Q(n491) );
  NAND4X0 U307 ( .IN1(n348), .IN2(instPacket_i[106]), .IN3(n342), .IN4(n340), 
        .QN(n434) );
  AOI22X1 U308 ( .IN1(n401), .IN2(n325), .IN3(n476), .IN4(n382), .QN(n431) );
  AO22X1 U309 ( .IN1(n351), .IN2(n354), .IN3(n444), .IN4(instPacket_i[103]), 
        .Q(n382) );
  NAND3X0 U310 ( .IN1(instPacket_i[103]), .IN2(n353), .IN3(instPacket_i[104]), 
        .QN(n436) );
  AOI222X1 U311 ( .IN1(n476), .IN2(n401), .IN3(n381), .IN4(n324), .IN5(n350), 
        .IN6(n325), .QN(n432) );
  NAND3X0 U312 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[101]), .IN3(n447), 
        .QN(n410) );
  AND3X1 U313 ( .IN1(instPacket_i[101]), .IN2(n353), .IN3(n447), .Q(n401) );
  AND2X1 U314 ( .IN1(n380), .IN2(instPacket_i[105]), .Q(n476) );
  AND3X1 U315 ( .IN1(n341), .IN2(n329), .IN3(instPacket_i[107]), .Q(n380) );
  AO21X1 U316 ( .IN1(n409), .IN2(n385), .IN3(n399), .Q(n384) );
  AND3X1 U317 ( .IN1(n396), .IN2(n404), .IN3(n397), .Q(n409) );
  AND2X1 U318 ( .IN1(n441), .IN2(n403), .Q(n397) );
  NAND3X0 U319 ( .IN1(instPacket_i[101]), .IN2(n379), .IN3(instPacket_i[102]), 
        .QN(n404) );
  NAND4X0 U320 ( .IN1(n331), .IN2(n406), .IN3(n378), .IN4(n455), .QN(n462) );
  NAND3X0 U321 ( .IN1(n379), .IN2(n353), .IN3(instPacket_i[101]), .QN(n385) );
  AND3X1 U322 ( .IN1(n353), .IN2(n352), .IN3(instPacket_i[104]), .Q(n375) );
  NAND3X0 U323 ( .IN1(n342), .IN2(n341), .IN3(n374), .QN(n399) );
  NOR3X0 U324 ( .IN1(n419), .IN2(n418), .IN3(n373), .QN(n406) );
  AOI21X1 U325 ( .IN1(n400), .IN2(n372), .IN3(n376), .QN(n373) );
  NAND3X0 U326 ( .IN1(n374), .IN2(n342), .IN3(instPacket_i[106]), .QN(n376) );
  NAND3X0 U327 ( .IN1(n379), .IN2(n354), .IN3(instPacket_i[102]), .QN(n396) );
  NAND3X0 U328 ( .IN1(n421), .IN2(n417), .IN3(n371), .QN(n425) );
  NAND3X0 U329 ( .IN1(n354), .IN2(n353), .IN3(n447), .QN(n372) );
  NAND3X0 U330 ( .IN1(instPacket_i[102]), .IN2(n354), .IN3(n447), .QN(n400) );
  AND3X1 U331 ( .IN1(instPacket_i[105]), .IN2(n374), .IN3(instPacket_i[106]), 
        .Q(n377) );
  NAND3X0 U332 ( .IN1(n354), .IN2(n353), .IN3(n379), .QN(n442) );
  HADDX1 \r339/U1_1_1  ( .A0(instPacket_i_86), .B0(instPacket_i_85), .C1(
        \r339/carry[2] ), .SO(N280) );
  HADDX1 \r339/U1_1_2  ( .A0(instPacket_i_87), .B0(\r339/carry[2] ), .C1(
        \r339/carry[3] ), .SO(N281) );
  HADDX1 \r339/U1_1_3  ( .A0(instPacket_i_88), .B0(\r339/carry[3] ), .C1(
        \r339/carry[4] ), .SO(N282) );
  HADDX1 \r339/U1_1_4  ( .A0(instPacket_i_89), .B0(\r339/carry[4] ), .C1(
        \r339/carry[5] ), .SO(N283) );
  INVX0 U3 ( .INP(1'b1), .ZN(decodedPacket1_o[5]) );
  INVX0 U5 ( .INP(1'b1), .ZN(decodedPacket1_o[6]) );
  INVX0 U7 ( .INP(1'b1), .ZN(decodedPacket1_o[7]) );
  INVX0 U9 ( .INP(1'b1), .ZN(decodedPacket1_o[8]) );
  INVX0 U11 ( .INP(1'b1), .ZN(decodedPacket1_o[9]) );
  INVX0 U13 ( .INP(1'b1), .ZN(decodedPacket1_o[10]) );
  INVX0 U15 ( .INP(1'b1), .ZN(decodedPacket1_o[11]) );
  INVX0 U17 ( .INP(1'b1), .ZN(decodedPacket1_o[12]) );
  INVX0 U19 ( .INP(1'b1), .ZN(decodedPacket1_o[13]) );
  INVX0 U21 ( .INP(1'b1), .ZN(decodedPacket1_o[14]) );
  INVX0 U23 ( .INP(1'b1), .ZN(decodedPacket1_o[15]) );
  INVX0 U25 ( .INP(1'b1), .ZN(decodedPacket1_o[16]) );
  INVX0 U27 ( .INP(1'b1), .ZN(decodedPacket1_o[17]) );
  INVX0 U29 ( .INP(1'b1), .ZN(decodedPacket1_o[18]) );
  INVX0 U31 ( .INP(1'b1), .ZN(decodedPacket1_o[19]) );
  INVX0 U33 ( .INP(1'b1), .ZN(decodedPacket1_o[20]) );
  INVX0 U35 ( .INP(1'b1), .ZN(decodedPacket1_o[21]) );
  INVX0 U37 ( .INP(1'b1), .ZN(decodedPacket1_o[22]) );
  INVX0 U39 ( .INP(1'b1), .ZN(decodedPacket1_o[23]) );
  INVX0 U41 ( .INP(1'b1), .ZN(decodedPacket1_o[24]) );
  INVX0 U43 ( .INP(1'b1), .ZN(decodedPacket1_o[25]) );
  INVX0 U45 ( .INP(1'b1), .ZN(decodedPacket1_o[26]) );
  INVX0 U47 ( .INP(1'b1), .ZN(decodedPacket1_o[27]) );
  INVX0 U49 ( .INP(1'b1), .ZN(decodedPacket1_o[28]) );
  INVX0 U51 ( .INP(1'b1), .ZN(decodedPacket1_o[29]) );
  INVX0 U53 ( .INP(1'b1), .ZN(decodedPacket1_o[30]) );
  INVX0 U55 ( .INP(1'b1), .ZN(decodedPacket1_o[31]) );
  INVX0 U57 ( .INP(1'b1), .ZN(decodedPacket1_o[32]) );
  INVX0 U59 ( .INP(1'b1), .ZN(decodedPacket1_o[33]) );
  INVX0 U61 ( .INP(1'b1), .ZN(decodedPacket1_o[34]) );
  INVX0 U63 ( .INP(1'b1), .ZN(decodedPacket1_o[35]) );
  INVX0 U65 ( .INP(1'b1), .ZN(decodedPacket1_o[36]) );
  INVX0 U67 ( .INP(1'b1), .ZN(decodedPacket1_o[117]) );
  INVX0 U69 ( .INP(1'b1), .ZN(decodedPacket1_o[121]) );
  INVX0 U71 ( .INP(1'b1), .ZN(decodedPacket1_o[122]) );
  INVX0 U73 ( .INP(1'b1), .ZN(decodedPacket1_o[123]) );
  INVX0 U75 ( .INP(1'b1), .ZN(decodedPacket1_o[124]) );
  INVX0 U77 ( .INP(1'b1), .ZN(decodedPacket1_o[125]) );
  INVX0 U79 ( .INP(1'b1), .ZN(decodedPacket0_o[122]) );
  INVX0 U81 ( .INP(1'b1), .ZN(decodedPacket0_o[123]) );
  INVX0 U83 ( .INP(1'b1), .ZN(decodedPacket0_o[124]) );
  INVX0 U85 ( .INP(1'b1), .ZN(decodedPacket0_o[125]) );
  INVX0 U87 ( .INP(decodedPacket1_o[77]), .ZN(n316) );
  NBUFFX2 U88 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[69]) );
  NBUFFX2 U89 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[73]) );
  NBUFFX2 U90 ( .INP(decodedPacket1_o[74]), .Z(decodedPacket1_o[75]) );
  NBUFFX2 U91 ( .INP(n511), .Z(decodedPacket1_o[74]) );
  NBUFFX2 U92 ( .INP(n511), .Z(decodedPacket1_o[77]) );
  NOR2X0 U93 ( .IN1(n506), .IN2(n459), .QN(n511) );
  INVX0 U94 ( .INP(n499), .ZN(n322) );
  NOR2X0 U95 ( .IN1(n336), .IN2(n308), .QN(decodedPacket1_o_119) );
  INVX0 U96 ( .INP(n482), .ZN(decodedPacket0_o[84]) );
  NBUFFX2 U97 ( .INP(n510), .Z(n314) );
  INVX0 U98 ( .INP(n509), .ZN(decodedPacket1_o[71]) );
  INVX0 U99 ( .INP(n468), .ZN(n317) );
  INVX0 U100 ( .INP(n500), .ZN(n318) );
  NOR2X0 U101 ( .IN1(n308), .IN2(n317), .QN(n472) );
  INVX0 U102 ( .INP(n460), .ZN(n321) );
  NAND2X1 U103 ( .IN1(n343), .IN2(n337), .QN(n489) );
  INVX0 U104 ( .INP(n423), .ZN(n334) );
  INVX0 U105 ( .INP(n485), .ZN(n323) );
  INVX0 U106 ( .INP(n412), .ZN(n338) );
  INVX0 U107 ( .INP(n467), .ZN(n319) );
  INVX0 U108 ( .INP(n463), .ZN(n320) );
  NOR2X0 U109 ( .IN1(n422), .IN2(n333), .QN(n455) );
  INVX0 U110 ( .INP(n424), .ZN(n333) );
  NAND2X1 U111 ( .IN1(n345), .IN2(n325), .QN(n456) );
  INVX0 U112 ( .INP(n478), .ZN(n326) );
  INVX0 U113 ( .INP(n443), .ZN(n325) );
  NOR2X0 U114 ( .IN1(n307), .IN2(n322), .QN(decodedPacket1_o[72]) );
  NAND2X1 U115 ( .IN1(n315), .IN2(n395), .QN(n402) );
  NAND2X1 U116 ( .IN1(n315), .IN2(n481), .QN(n482) );
  INVX0 U117 ( .INP(n506), .ZN(n315) );
  NOR2X0 U118 ( .IN1(n412), .IN2(n405), .QN(n378) );
  NOR2X0 U119 ( .IN1(n308), .IN2(n455), .QN(decodedPacket1_o_118) );
  NOR4X0 U120 ( .IN1(n464), .IN2(n463), .IN3(n478), .IN4(n462), .QN(n465) );
  NOR2X0 U121 ( .IN1(n307), .IN2(n424), .QN(decodedPacket1_o_120) );
  INVX0 U122 ( .INP(n399), .ZN(n337) );
  INVX0 U123 ( .INP(n442), .ZN(n343) );
  NOR2X0 U124 ( .IN1(n440), .IN2(n399), .QN(n412) );
  NOR2X0 U125 ( .IN1(n420), .IN2(n307), .QN(decodedPacket0_o[117]) );
  INVX0 U126 ( .INP(n417), .ZN(n332) );
  NOR2X0 U127 ( .IN1(n416), .IN2(n307), .QN(decodedPacket0_o[116]) );
  NOR4X0 U128 ( .IN1(n415), .IN2(n414), .IN3(n425), .IN4(n423), .QN(n416) );
  NOR2X0 U129 ( .IN1(n487), .IN2(n307), .QN(decodedPacket0_o[91]) );
  NOR4X0 U130 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(n487) );
  OR2X1 U131 ( .IN1(decodedPacket1_o[118]), .IN2(n224), .Q(
        decodedPacket0_o[118]) );
  AOI21X1 U132 ( .IN1(n335), .IN2(n421), .IN3(n308), .QN(n224) );
  INVX0 U133 ( .INP(n372), .ZN(n349) );
  INVX0 U134 ( .INP(n422), .ZN(n336) );
  NOR2X0 U135 ( .IN1(n474), .IN2(n308), .QN(n471) );
  NOR2X0 U136 ( .IN1(n343), .IN2(n346), .QN(n426) );
  OA21X1 U137 ( .IN1(n395), .IN2(n328), .IN3(n315), .Q(decodedPacket0_o[98])
         );
  INVX0 U138 ( .INP(n474), .ZN(n328) );
  NAND2X1 U139 ( .IN1(n406), .IN2(n335), .QN(n423) );
  INVX0 U140 ( .INP(n405), .ZN(n335) );
  INVX0 U141 ( .INP(n492), .ZN(n339) );
  NAND2X1 U142 ( .IN1(n315), .IN2(n457), .QN(n509) );
  NOR2X0 U143 ( .IN1(n350), .IN2(n345), .QN(n428) );
  INVX0 U144 ( .INP(n425), .ZN(n331) );
  NAND2X1 U145 ( .IN1(n473), .IN2(n474), .QN(n467) );
  INVX0 U146 ( .INP(n484), .ZN(n327) );
  INVX0 U147 ( .INP(n396), .ZN(n345) );
  NOR2X0 U148 ( .IN1(n403), .IN2(n376), .QN(n422) );
  INVX0 U149 ( .INP(n385), .ZN(n346) );
  NOR2X0 U150 ( .IN1(n443), .IN2(n403), .QN(n478) );
  NAND2X1 U151 ( .IN1(n346), .IN2(n377), .QN(n424) );
  NAND2X1 U152 ( .IN1(n380), .IN2(n342), .QN(n443) );
  NAND2X1 U153 ( .IN1(n375), .IN2(n354), .QN(n441) );
  INVX0 U154 ( .INP(n462), .ZN(n330) );
  NAND2X1 U155 ( .IN1(n349), .IN2(n377), .QN(n371) );
  NOR2X0 U156 ( .IN1(n441), .IN2(n376), .QN(n405) );
  NOR2X0 U157 ( .IN1(n442), .IN2(n376), .QN(n418) );
  NOR2X0 U158 ( .IN1(n396), .IN2(n376), .QN(n419) );
  NOR2X0 U159 ( .IN1(n400), .IN2(n399), .QN(n492) );
  NOR2X0 U274 ( .IN1(n370), .IN2(n402), .QN(decodedPacket0_o[107]) );
  NOR2X0 U298 ( .IN1(n369), .IN2(n402), .QN(decodedPacket0_o[108]) );
  NOR2X0 U333 ( .IN1(n368), .IN2(n402), .QN(decodedPacket0_o[109]) );
  NOR2X0 U334 ( .IN1(n367), .IN2(n402), .QN(decodedPacket0_o[110]) );
  NOR2X0 U335 ( .IN1(n366), .IN2(n402), .QN(decodedPacket0_o[111]) );
  NAND2X1 U336 ( .IN1(n476), .IN2(n386), .QN(n474) );
  NOR2X0 U337 ( .IN1(n362), .IN2(n482), .QN(decodedPacket0_o[85]) );
  NOR2X0 U338 ( .IN1(n361), .IN2(n482), .QN(decodedPacket0_o[86]) );
  NOR2X0 U339 ( .IN1(n360), .IN2(n482), .QN(decodedPacket0_o[87]) );
  NOR2X0 U340 ( .IN1(n359), .IN2(n482), .QN(decodedPacket0_o[88]) );
  NOR2X0 U341 ( .IN1(n358), .IN2(n482), .QN(decodedPacket0_o[89]) );
  NOR2X0 U342 ( .IN1(n357), .IN2(n482), .QN(decodedPacket0_o[90]) );
  NAND2X1 U343 ( .IN1(n316), .IN2(n342), .QN(decodedPacket0_o[73]) );
  NAND2X1 U344 ( .IN1(n316), .IN2(n341), .QN(decodedPacket0_o[74]) );
  NAND2X1 U345 ( .IN1(n316), .IN2(n340), .QN(decodedPacket0_o[75]) );
  NAND2X1 U346 ( .IN1(n316), .IN2(n329), .QN(decodedPacket0_o[76]) );
  NOR2X0 U347 ( .IN1(n475), .IN2(n308), .QN(decodedPacket0_o[83]) );
  NOR2X0 U348 ( .IN1(n496), .IN2(n307), .QN(decodedPacket0_o[94]) );
  NOR2X0 U349 ( .IN1(n497), .IN2(n308), .QN(decodedPacket0_o[95]) );
  NOR2X0 U350 ( .IN1(n494), .IN2(n308), .QN(decodedPacket0_o[92]) );
  NOR2X0 U351 ( .IN1(n492), .IN2(n503), .QN(n493) );
  NOR2X0 U352 ( .IN1(n498), .IN2(n307), .QN(decodedPacket0_o[96]) );
  NOR2X0 U353 ( .IN1(n470), .IN2(n308), .QN(decodedPacket0_o[78]) );
  NOR2X0 U354 ( .IN1(n495), .IN2(n308), .QN(decodedPacket0_o[93]) );
  INVX0 U355 ( .INP(n400), .ZN(n348) );
  NAND2X1 U356 ( .IN1(n509), .IN2(n352), .QN(decodedPacket0_o[71]) );
  NOR2X0 U357 ( .IN1(n436), .IN2(n427), .QN(n502) );
  INVX0 U358 ( .INP(n410), .ZN(n350) );
  NOR2X0 U359 ( .IN1(n316), .IN2(n356), .QN(decodedPacket1_o[78]) );
  NOR2X0 U360 ( .IN1(n316), .IN2(n355), .QN(decodedPacket1_o[83]) );
  NOR2X0 U361 ( .IN1(n352), .IN2(n443), .QN(n445) );
  NAND2X1 U362 ( .IN1(n444), .IN2(n352), .QN(n440) );
  NAND2X1 U363 ( .IN1(n348), .IN2(n377), .QN(n417) );
  NAND2X1 U364 ( .IN1(n343), .IN2(n377), .QN(n421) );
  NAND2X1 U365 ( .IN1(n476), .IN2(n344), .QN(n429) );
  NOR2X0 U366 ( .IN1(n503), .IN2(n502), .QN(n430) );
  INVX0 U367 ( .INP(n428), .ZN(n344) );
  NOR2X0 U368 ( .IN1(n501), .IN2(n357), .QN(n504) );
  NAND2X1 U369 ( .IN1(n350), .IN2(n476), .QN(n383) );
  NAND2X1 U370 ( .IN1(n476), .IN2(n345), .QN(n477) );
  INVX0 U371 ( .INP(n436), .ZN(n351) );
  NAND2X1 U372 ( .IN1(n337), .IN2(n411), .QN(n413) );
  INVX0 U373 ( .INP(n427), .ZN(n324) );
  NOR2X0 U374 ( .IN1(n352), .IN2(n450), .QN(n381) );
  NBUFFX2 U375 ( .INP(instPacketValid_i), .Z(decodedPacket0Valid_o) );
  NOR2X0 U376 ( .IN1(n352), .IN2(instPacket_i[104]), .QN(n379) );
  NAND2X1 U377 ( .IN1(n375), .IN2(instPacket_i[101]), .QN(n403) );
  INVX0 U378 ( .INP(instPacket_i[103]), .ZN(n352) );
  INVX0 U379 ( .INP(instPacket_i[101]), .ZN(n354) );
  INVX0 U380 ( .INP(instPacket_i[105]), .ZN(n342) );
  INVX0 U381 ( .INP(instPacket_i[102]), .ZN(n353) );
  INVX0 U382 ( .INP(instPacket_i[106]), .ZN(n341) );
  NOR2X0 U383 ( .IN1(instPacket_i[108]), .IN2(instPacket_i[107]), .QN(n374) );
  INVX0 U384 ( .INP(instPacket_i[108]), .ZN(n329) );
  NOR4X0 U385 ( .IN1(n390), .IN2(instPacket_i[127]), .IN3(instPacket_i[129]), 
        .IN4(instPacket_i[128]), .QN(n391) );
  NOR4X0 U386 ( .IN1(n389), .IN2(instPacket_i[121]), .IN3(instPacket_i[123]), 
        .IN4(instPacket_i[122]), .QN(n392) );
  NOR4X0 U387 ( .IN1(n387), .IN2(instPacket_i[109]), .IN3(instPacket_i[111]), 
        .IN4(instPacket_i[110]), .QN(n394) );
  NOR4X0 U388 ( .IN1(n388), .IN2(instPacket_i[115]), .IN3(instPacket_i[117]), 
        .IN4(instPacket_i[116]), .QN(n393) );
  NOR4X0 U389 ( .IN1(n483), .IN2(n484), .IN3(n307), .IN4(n452), .QN(n453) );
  NOR2X0 U390 ( .IN1(n365), .IN2(n402), .QN(decodedPacket0_o[112]) );
  INVX0 U391 ( .INP(instPacket_i_82), .ZN(n365) );
  NOR2X0 U392 ( .IN1(n364), .IN2(n402), .QN(decodedPacket0_o[113]) );
  INVX0 U393 ( .INP(instPacket_i_83), .ZN(n364) );
  NOR2X0 U394 ( .IN1(n363), .IN2(n402), .QN(decodedPacket0_o[114]) );
  INVX0 U395 ( .INP(instPacket_i_84), .ZN(n363) );
  INVX0 U396 ( .INP(n447), .ZN(n347) );
  NOR2X0 U397 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[102]), .QN(n448) );
  NOR2X0 U398 ( .IN1(n507), .IN2(n307), .QN(decodedPacket0_o[97]) );
  NOR4X0 U399 ( .IN1(n505), .IN2(n504), .IN3(n503), .IN4(n502), .QN(n507) );
  NOR2X0 U400 ( .IN1(instPacket_i[104]), .IN2(instPacket_i[103]), .QN(n447) );
  NBUFFX2 U401 ( .INP(instPacket_i[45]), .Z(decodedPacket0_o[45]) );
  NBUFFX2 U402 ( .INP(instPacket_i[46]), .Z(decodedPacket0_o[46]) );
  NBUFFX2 U403 ( .INP(instPacket_i[47]), .Z(decodedPacket0_o[47]) );
  NBUFFX2 U404 ( .INP(instPacket_i[48]), .Z(decodedPacket0_o[48]) );
  NBUFFX2 U405 ( .INP(instPacket_i[49]), .Z(decodedPacket0_o[49]) );
  NBUFFX2 U406 ( .INP(instPacket_i[50]), .Z(decodedPacket0_o[50]) );
  NBUFFX2 U407 ( .INP(instPacket_i[51]), .Z(decodedPacket0_o[51]) );
  NBUFFX2 U408 ( .INP(instPacket_i[52]), .Z(decodedPacket0_o[52]) );
  NBUFFX2 U409 ( .INP(instPacket_i[53]), .Z(decodedPacket0_o[53]) );
  NBUFFX2 U410 ( .INP(instPacket_i[54]), .Z(decodedPacket0_o[54]) );
  NBUFFX2 U411 ( .INP(instPacket_i[55]), .Z(decodedPacket0_o[55]) );
  NBUFFX2 U412 ( .INP(instPacket_i[56]), .Z(decodedPacket0_o[56]) );
  NBUFFX2 U413 ( .INP(instPacket_i[57]), .Z(decodedPacket0_o[57]) );
  NBUFFX2 U414 ( .INP(instPacket_i[58]), .Z(decodedPacket0_o[58]) );
  NBUFFX2 U415 ( .INP(instPacket_i[59]), .Z(decodedPacket0_o[59]) );
  NBUFFX2 U416 ( .INP(instPacket_i[60]), .Z(decodedPacket0_o[60]) );
  NBUFFX2 U417 ( .INP(instPacket_i[61]), .Z(decodedPacket0_o[61]) );
  NBUFFX2 U418 ( .INP(instPacket_i[62]), .Z(decodedPacket0_o[62]) );
  NBUFFX2 U419 ( .INP(instPacket_i[63]), .Z(decodedPacket0_o[63]) );
  NBUFFX2 U420 ( .INP(instPacket_i[64]), .Z(decodedPacket0_o[64]) );
  NBUFFX2 U421 ( .INP(instPacket_i[65]), .Z(decodedPacket0_o[65]) );
  NBUFFX2 U422 ( .INP(instPacket_i[66]), .Z(decodedPacket0_o[66]) );
  NBUFFX2 U423 ( .INP(instPacket_i[67]), .Z(decodedPacket0_o[67]) );
  NBUFFX2 U424 ( .INP(instPacket_i[68]), .Z(decodedPacket0_o[68]) );
  NAND2X1 U425 ( .IN1(instPacket_i[102]), .IN2(instPacket_i[104]), .QN(n450)
         );
  NOR2X0 U426 ( .IN1(n450), .IN2(instPacket_i[101]), .QN(n444) );
  INVX0 U427 ( .INP(instPacket_i_71), .ZN(N287) );
  XNOR2X1 U428 ( .IN1(n225), .IN2(instPacket_i_84), .Q(N300) );
  NAND2X1 U429 ( .IN1(instPacket_i_83), .IN2(\r340/carry[14] ), .QN(n225) );
  NBUFFX2 U430 ( .INP(instPacket_i[45]), .Z(decodedPacket1_o[45]) );
  NBUFFX2 U431 ( .INP(instPacket_i[46]), .Z(decodedPacket1_o[46]) );
  NBUFFX2 U432 ( .INP(instPacket_i[47]), .Z(decodedPacket1_o[47]) );
  NBUFFX2 U433 ( .INP(instPacket_i[48]), .Z(decodedPacket1_o[48]) );
  NBUFFX2 U434 ( .INP(instPacket_i[49]), .Z(decodedPacket1_o[49]) );
  NBUFFX2 U435 ( .INP(instPacket_i[50]), .Z(decodedPacket1_o[50]) );
  NBUFFX2 U436 ( .INP(instPacket_i[51]), .Z(decodedPacket1_o[51]) );
  NBUFFX2 U437 ( .INP(instPacket_i[52]), .Z(decodedPacket1_o[52]) );
  NBUFFX2 U438 ( .INP(instPacket_i[53]), .Z(decodedPacket1_o[53]) );
  NBUFFX2 U439 ( .INP(instPacket_i[54]), .Z(decodedPacket1_o[54]) );
  NBUFFX2 U440 ( .INP(instPacket_i[55]), .Z(decodedPacket1_o[55]) );
  NBUFFX2 U441 ( .INP(instPacket_i[56]), .Z(decodedPacket1_o[56]) );
  NBUFFX2 U442 ( .INP(instPacket_i[57]), .Z(decodedPacket1_o[57]) );
  NBUFFX2 U443 ( .INP(instPacket_i[58]), .Z(decodedPacket1_o[58]) );
  NBUFFX2 U444 ( .INP(instPacket_i[59]), .Z(decodedPacket1_o[59]) );
  NBUFFX2 U445 ( .INP(instPacket_i[60]), .Z(decodedPacket1_o[60]) );
  NBUFFX2 U446 ( .INP(instPacket_i[61]), .Z(decodedPacket1_o[61]) );
  NBUFFX2 U447 ( .INP(instPacket_i[62]), .Z(decodedPacket1_o[62]) );
  NBUFFX2 U448 ( .INP(instPacket_i[63]), .Z(decodedPacket1_o[63]) );
  NBUFFX2 U449 ( .INP(instPacket_i[64]), .Z(decodedPacket1_o[64]) );
  NBUFFX2 U450 ( .INP(instPacket_i[65]), .Z(decodedPacket1_o[65]) );
  NBUFFX2 U451 ( .INP(instPacket_i[66]), .Z(decodedPacket1_o[66]) );
  NBUFFX2 U452 ( .INP(instPacket_i[67]), .Z(decodedPacket1_o[67]) );
  NBUFFX2 U453 ( .INP(instPacket_i[68]), .Z(decodedPacket1_o[68]) );
  INVX0 U454 ( .INP(instPacket_i[107]), .ZN(n340) );
  INVX0 U455 ( .INP(instPacket_i_90), .ZN(n357) );
  NAND2X1 U456 ( .IN1(n325), .IN2(instPacket_i[101]), .QN(n427) );
  NOR2X0 U457 ( .IN1(n437), .IN2(n354), .QN(n438) );
  INVX0 U458 ( .INP(instPacket_i_85), .ZN(n362) );
  INVX0 U459 ( .INP(instPacket_i_93), .ZN(n356) );
  INVX0 U460 ( .INP(instPacket_i_98), .ZN(n355) );
  INVX0 U461 ( .INP(instPacket_i_77), .ZN(n370) );
  INVX0 U462 ( .INP(instPacket_i_78), .ZN(n369) );
  INVX0 U463 ( .INP(instPacket_i_79), .ZN(n368) );
  INVX0 U464 ( .INP(instPacket_i_80), .ZN(n367) );
  INVX0 U465 ( .INP(instPacket_i_81), .ZN(n366) );
  INVX0 U466 ( .INP(instPacket_i_86), .ZN(n361) );
  INVX0 U467 ( .INP(instPacket_i_87), .ZN(n360) );
  INVX0 U468 ( .INP(instPacket_i_88), .ZN(n359) );
  INVX0 U469 ( .INP(instPacket_i_89), .ZN(n358) );
  NBUFFX2 U470 ( .INP(instPacket_i[44]), .Z(decodedPacket0_o[44]) );
  NBUFFX2 U471 ( .INP(instPacket_i[44]), .Z(decodedPacket1_o[44]) );
  NBUFFX2 U472 ( .INP(instPacket_i[43]), .Z(decodedPacket0_o[43]) );
  NBUFFX2 U473 ( .INP(instPacket_i[43]), .Z(decodedPacket1_o[43]) );
  NBUFFX2 U474 ( .INP(instPacket_i[42]), .Z(decodedPacket0_o[42]) );
  NBUFFX2 U475 ( .INP(instPacket_i[42]), .Z(decodedPacket1_o[42]) );
  NBUFFX2 U476 ( .INP(instPacket_i[41]), .Z(decodedPacket0_o[41]) );
  NBUFFX2 U477 ( .INP(instPacket_i[41]), .Z(decodedPacket1_o[41]) );
  NBUFFX2 U478 ( .INP(instPacket_i[40]), .Z(decodedPacket0_o[40]) );
  NBUFFX2 U479 ( .INP(instPacket_i[40]), .Z(decodedPacket1_o[40]) );
  NBUFFX2 U480 ( .INP(instPacket_i[39]), .Z(decodedPacket0_o[39]) );
  NBUFFX2 U481 ( .INP(instPacket_i[39]), .Z(decodedPacket1_o[39]) );
  NBUFFX2 U482 ( .INP(instPacket_i[38]), .Z(decodedPacket0_o[38]) );
  NBUFFX2 U483 ( .INP(instPacket_i[38]), .Z(decodedPacket1_o[38]) );
  NBUFFX2 U484 ( .INP(instPacket_i[37]), .Z(decodedPacket0_o[37]) );
  NBUFFX2 U485 ( .INP(instPacket_i[37]), .Z(decodedPacket1_o[37]) );
  NBUFFX2 U486 ( .INP(instPacket_i[4]), .Z(decodedPacket0_o[4]) );
  NBUFFX2 U487 ( .INP(instPacket_i[4]), .Z(decodedPacket1_o[4]) );
  NBUFFX2 U488 ( .INP(instPacket_i[3]), .Z(decodedPacket0_o[3]) );
  NBUFFX2 U489 ( .INP(instPacket_i[3]), .Z(decodedPacket1_o[3]) );
  NBUFFX2 U490 ( .INP(instPacket_i[2]), .Z(decodedPacket0_o[2]) );
  NBUFFX2 U491 ( .INP(instPacket_i[2]), .Z(decodedPacket1_o[2]) );
  NBUFFX2 U492 ( .INP(instPacket_i[1]), .Z(decodedPacket0_o[1]) );
  NBUFFX2 U493 ( .INP(instPacket_i[1]), .Z(decodedPacket1_o[1]) );
  NBUFFX2 U494 ( .INP(instPacket_i[0]), .Z(decodedPacket0_o[0]) );
  NBUFFX2 U495 ( .INP(instPacket_i[0]), .Z(decodedPacket1_o[0]) );
  NBUFFX2 U496 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[98]) );
  NBUFFX2 U497 ( .INP(decodedPacket1_o_118), .Z(decodedPacket1_o[118]) );
  NBUFFX2 U498 ( .INP(decodedPacket1_o[76]), .Z(decodedPacket1_o[115]) );
  NBUFFX2 U499 ( .INP(n511), .Z(decodedPacket1_o[76]) );
  NBUFFX2 U500 ( .INP(n508), .Z(n312) );
  NBUFFX2 U501 ( .INP(n510), .Z(decodedPacket0_o[121]) );
  NAND4X0 U502 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n307) );
  NAND4X0 U503 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n308) );
  XOR2X1 U504 ( .IN1(\r340/carry[14] ), .IN2(instPacket_i_83), .Q(N299) );
  AND2X1 U505 ( .IN1(instPacket_i_82), .IN2(\r340/carry[13] ), .Q(
        \r340/carry[14] ) );
  XOR2X1 U506 ( .IN1(\r340/carry[13] ), .IN2(instPacket_i_82), .Q(N298) );
  AND2X1 U507 ( .IN1(instPacket_i_81), .IN2(\r340/carry[12] ), .Q(
        \r340/carry[13] ) );
  XOR2X1 U508 ( .IN1(\r340/carry[12] ), .IN2(instPacket_i_81), .Q(N297) );
  AND2X1 U509 ( .IN1(instPacket_i_80), .IN2(\r340/carry[11] ), .Q(
        \r340/carry[12] ) );
  XOR2X1 U510 ( .IN1(\r340/carry[11] ), .IN2(instPacket_i_80), .Q(N296) );
  AND2X1 U511 ( .IN1(instPacket_i_79), .IN2(\r340/carry[10] ), .Q(
        \r340/carry[11] ) );
  XOR2X1 U512 ( .IN1(\r340/carry[10] ), .IN2(instPacket_i_79), .Q(N295) );
  AND2X1 U513 ( .IN1(instPacket_i_78), .IN2(\r340/carry[9] ), .Q(
        \r340/carry[10] ) );
  XOR2X1 U514 ( .IN1(\r340/carry[9] ), .IN2(instPacket_i_78), .Q(N294) );
  AND2X1 U515 ( .IN1(instPacket_i_77), .IN2(\r340/carry[8] ), .Q(
        \r340/carry[9] ) );
  XOR2X1 U516 ( .IN1(\r340/carry[8] ), .IN2(instPacket_i_77), .Q(N293) );
  AND2X1 U517 ( .IN1(instPacket_i_76), .IN2(\r340/carry[7] ), .Q(
        \r340/carry[8] ) );
  XOR2X1 U518 ( .IN1(\r340/carry[7] ), .IN2(instPacket_i_76), .Q(N292) );
  AND2X1 U519 ( .IN1(instPacket_i_75), .IN2(\r340/carry[6] ), .Q(
        \r340/carry[7] ) );
  XOR2X1 U520 ( .IN1(\r340/carry[6] ), .IN2(instPacket_i_75), .Q(N291) );
  AND2X1 U521 ( .IN1(instPacket_i_74), .IN2(\r340/carry[5] ), .Q(
        \r340/carry[6] ) );
  XOR2X1 U522 ( .IN1(\r340/carry[5] ), .IN2(instPacket_i_74), .Q(N290) );
  AND2X1 U523 ( .IN1(instPacket_i_73), .IN2(\r340/carry[4] ), .Q(
        \r340/carry[5] ) );
  XOR2X1 U524 ( .IN1(\r340/carry[4] ), .IN2(instPacket_i_73), .Q(N289) );
  AND2X1 U525 ( .IN1(instPacket_i_72), .IN2(instPacket_i_71), .Q(
        \r340/carry[4] ) );
  XOR2X1 U526 ( .IN1(instPacket_i_71), .IN2(instPacket_i_72), .Q(N288) );
  XOR2X1 U527 ( .IN1(\r339/carry[5] ), .IN2(instPacket_i_90), .Q(N284) );
endmodule


module Decode ( reset, clk, fs2Ready_i, inst0PacketValid_i, inst0Packet_i, 
        inst1PacketValid_i, inst1Packet_i, inst2PacketValid_i, inst2Packet_i, 
        inst3PacketValid_i, inst3Packet_i, decodeReady_o, decodedVector_o, 
        decodedPacket0_o, decodedPacket1_o, decodedPacket2_o, decodedPacket3_o, 
        decodedPacket4_o, decodedPacket5_o, decodedPacket6_o, decodedPacket7_o
 );
  input [132:0] inst0Packet_i;
  input [132:0] inst1Packet_i;
  input [132:0] inst2Packet_i;
  input [132:0] inst3Packet_i;
  output [7:0] decodedVector_o;
  output [125:0] decodedPacket0_o;
  output [125:0] decodedPacket1_o;
  output [125:0] decodedPacket2_o;
  output [125:0] decodedPacket3_o;
  output [125:0] decodedPacket4_o;
  output [125:0] decodedPacket5_o;
  output [125:0] decodedPacket6_o;
  output [125:0] decodedPacket7_o;
  input reset, clk, fs2Ready_i, inst0PacketValid_i, inst1PacketValid_i,
         inst2PacketValid_i, inst3PacketValid_i;
  output decodeReady_o;
  wire   \decodedPacket[7][120] , \decodedPacket[7][119] ,
         \decodedPacket[7][118] , \decodedPacket[7][116] ,
         \decodedPacket[7][115] , \decodedPacket[7][114] ,
         \decodedPacket[7][113] , \decodedPacket[7][112] ,
         \decodedPacket[7][111] , \decodedPacket[7][110] ,
         \decodedPacket[7][109] , \decodedPacket[7][108] ,
         \decodedPacket[7][107] , \decodedPacket[7][106] ,
         \decodedPacket[7][105] , \decodedPacket[7][104] ,
         \decodedPacket[7][103] , \decodedPacket[7][102] ,
         \decodedPacket[7][101] , \decodedPacket[7][100] ,
         \decodedPacket[7][99] , \decodedPacket[7][98] ,
         \decodedPacket[7][97] , \decodedPacket[7][96] ,
         \decodedPacket[7][95] , \decodedPacket[7][94] ,
         \decodedPacket[7][93] , \decodedPacket[7][92] ,
         \decodedPacket[7][91] , \decodedPacket[7][90] ,
         \decodedPacket[7][89] , \decodedPacket[7][88] ,
         \decodedPacket[7][87] , \decodedPacket[7][86] ,
         \decodedPacket[7][85] , \decodedPacket[7][84] ,
         \decodedPacket[7][83] , \decodedPacket[7][82] ,
         \decodedPacket[7][81] , \decodedPacket[7][80] ,
         \decodedPacket[7][79] , \decodedPacket[7][78] ,
         \decodedPacket[7][77] , \decodedPacket[7][76] ,
         \decodedPacket[7][75] , \decodedPacket[7][74] ,
         \decodedPacket[7][73] , \decodedPacket[7][72] ,
         \decodedPacket[7][71] , \decodedPacket[7][70] ,
         \decodedPacket[7][69] , \decodedPacket[7][68] ,
         \decodedPacket[7][67] , \decodedPacket[7][66] ,
         \decodedPacket[7][65] , \decodedPacket[7][64] ,
         \decodedPacket[7][63] , \decodedPacket[7][62] ,
         \decodedPacket[7][61] , \decodedPacket[7][60] ,
         \decodedPacket[7][59] , \decodedPacket[7][58] ,
         \decodedPacket[7][57] , \decodedPacket[7][56] ,
         \decodedPacket[7][55] , \decodedPacket[7][54] ,
         \decodedPacket[7][53] , \decodedPacket[7][52] ,
         \decodedPacket[7][51] , \decodedPacket[7][50] ,
         \decodedPacket[7][49] , \decodedPacket[7][48] ,
         \decodedPacket[7][47] , \decodedPacket[7][46] ,
         \decodedPacket[7][45] , \decodedPacket[7][44] ,
         \decodedPacket[7][43] , \decodedPacket[7][42] ,
         \decodedPacket[7][41] , \decodedPacket[7][40] ,
         \decodedPacket[7][39] , \decodedPacket[7][38] ,
         \decodedPacket[7][37] , \decodedPacket[7][4] , \decodedPacket[7][3] ,
         \decodedPacket[7][2] , \decodedPacket[7][1] , \decodedPacket[7][0] ,
         \decodedPacket[6][121] , \decodedPacket[6][120] ,
         \decodedPacket[6][119] , \decodedPacket[6][118] ,
         \decodedPacket[6][117] , \decodedPacket[6][116] ,
         \decodedPacket[6][115] , \decodedPacket[6][114] ,
         \decodedPacket[6][113] , \decodedPacket[6][112] ,
         \decodedPacket[6][111] , \decodedPacket[6][110] ,
         \decodedPacket[6][109] , \decodedPacket[6][108] ,
         \decodedPacket[6][107] , \decodedPacket[6][106] ,
         \decodedPacket[6][105] , \decodedPacket[6][104] ,
         \decodedPacket[6][103] , \decodedPacket[6][102] ,
         \decodedPacket[6][101] , \decodedPacket[6][100] ,
         \decodedPacket[6][99] , \decodedPacket[6][98] ,
         \decodedPacket[6][97] , \decodedPacket[6][96] ,
         \decodedPacket[6][95] , \decodedPacket[6][94] ,
         \decodedPacket[6][93] , \decodedPacket[6][92] ,
         \decodedPacket[6][91] , \decodedPacket[6][90] ,
         \decodedPacket[6][89] , \decodedPacket[6][88] ,
         \decodedPacket[6][87] , \decodedPacket[6][86] ,
         \decodedPacket[6][85] , \decodedPacket[6][84] ,
         \decodedPacket[6][83] , \decodedPacket[6][82] ,
         \decodedPacket[6][81] , \decodedPacket[6][80] ,
         \decodedPacket[6][79] , \decodedPacket[6][78] ,
         \decodedPacket[6][77] , \decodedPacket[6][76] ,
         \decodedPacket[6][75] , \decodedPacket[6][74] ,
         \decodedPacket[6][73] , \decodedPacket[6][72] ,
         \decodedPacket[6][71] , \decodedPacket[6][70] ,
         \decodedPacket[6][69] , \decodedPacket[6][68] ,
         \decodedPacket[6][67] , \decodedPacket[6][66] ,
         \decodedPacket[6][65] , \decodedPacket[6][64] ,
         \decodedPacket[6][63] , \decodedPacket[6][62] ,
         \decodedPacket[6][61] , \decodedPacket[6][60] ,
         \decodedPacket[6][59] , \decodedPacket[6][58] ,
         \decodedPacket[6][57] , \decodedPacket[6][56] ,
         \decodedPacket[6][55] , \decodedPacket[6][54] ,
         \decodedPacket[6][53] , \decodedPacket[6][52] ,
         \decodedPacket[6][51] , \decodedPacket[6][50] ,
         \decodedPacket[6][49] , \decodedPacket[6][48] ,
         \decodedPacket[6][47] , \decodedPacket[6][46] ,
         \decodedPacket[6][45] , \decodedPacket[6][44] ,
         \decodedPacket[6][43] , \decodedPacket[6][42] ,
         \decodedPacket[6][41] , \decodedPacket[6][40] ,
         \decodedPacket[6][39] , \decodedPacket[6][38] ,
         \decodedPacket[6][37] , \decodedPacket[6][36] ,
         \decodedPacket[6][35] , \decodedPacket[6][34] ,
         \decodedPacket[6][33] , \decodedPacket[6][32] ,
         \decodedPacket[6][31] , \decodedPacket[6][30] ,
         \decodedPacket[6][29] , \decodedPacket[6][28] ,
         \decodedPacket[6][27] , \decodedPacket[6][26] ,
         \decodedPacket[6][25] , \decodedPacket[6][24] ,
         \decodedPacket[6][23] , \decodedPacket[6][22] ,
         \decodedPacket[6][21] , \decodedPacket[6][20] ,
         \decodedPacket[6][19] , \decodedPacket[6][18] ,
         \decodedPacket[6][17] , \decodedPacket[6][16] ,
         \decodedPacket[6][15] , \decodedPacket[6][14] ,
         \decodedPacket[6][13] , \decodedPacket[6][12] ,
         \decodedPacket[6][11] , \decodedPacket[6][10] , \decodedPacket[6][9] ,
         \decodedPacket[6][8] , \decodedPacket[6][7] , \decodedPacket[6][6] ,
         \decodedPacket[6][5] , \decodedPacket[6][4] , \decodedPacket[6][3] ,
         \decodedPacket[6][2] , \decodedPacket[6][1] , \decodedPacket[6][0] ,
         \decodedPacket[5][120] , \decodedPacket[5][119] ,
         \decodedPacket[5][118] , \decodedPacket[5][116] ,
         \decodedPacket[5][115] , \decodedPacket[5][114] ,
         \decodedPacket[5][113] , \decodedPacket[5][112] ,
         \decodedPacket[5][111] , \decodedPacket[5][110] ,
         \decodedPacket[5][109] , \decodedPacket[5][108] ,
         \decodedPacket[5][107] , \decodedPacket[5][106] ,
         \decodedPacket[5][105] , \decodedPacket[5][104] ,
         \decodedPacket[5][103] , \decodedPacket[5][102] ,
         \decodedPacket[5][101] , \decodedPacket[5][100] ,
         \decodedPacket[5][99] , \decodedPacket[5][98] ,
         \decodedPacket[5][97] , \decodedPacket[5][96] ,
         \decodedPacket[5][95] , \decodedPacket[5][94] ,
         \decodedPacket[5][93] , \decodedPacket[5][92] ,
         \decodedPacket[5][91] , \decodedPacket[5][90] ,
         \decodedPacket[5][89] , \decodedPacket[5][88] ,
         \decodedPacket[5][87] , \decodedPacket[5][86] ,
         \decodedPacket[5][85] , \decodedPacket[5][84] ,
         \decodedPacket[5][83] , \decodedPacket[5][82] ,
         \decodedPacket[5][81] , \decodedPacket[5][80] ,
         \decodedPacket[5][79] , \decodedPacket[5][78] ,
         \decodedPacket[5][77] , \decodedPacket[5][76] ,
         \decodedPacket[5][75] , \decodedPacket[5][74] ,
         \decodedPacket[5][73] , \decodedPacket[5][72] ,
         \decodedPacket[5][71] , \decodedPacket[5][70] ,
         \decodedPacket[5][69] , \decodedPacket[5][68] ,
         \decodedPacket[5][67] , \decodedPacket[5][66] ,
         \decodedPacket[5][65] , \decodedPacket[5][64] ,
         \decodedPacket[5][63] , \decodedPacket[5][62] ,
         \decodedPacket[5][61] , \decodedPacket[5][60] ,
         \decodedPacket[5][59] , \decodedPacket[5][58] ,
         \decodedPacket[5][57] , \decodedPacket[5][56] ,
         \decodedPacket[5][55] , \decodedPacket[5][54] ,
         \decodedPacket[5][53] , \decodedPacket[5][52] ,
         \decodedPacket[5][51] , \decodedPacket[5][50] ,
         \decodedPacket[5][49] , \decodedPacket[5][48] ,
         \decodedPacket[5][47] , \decodedPacket[5][46] ,
         \decodedPacket[5][45] , \decodedPacket[5][44] ,
         \decodedPacket[5][43] , \decodedPacket[5][42] ,
         \decodedPacket[5][41] , \decodedPacket[5][40] ,
         \decodedPacket[5][39] , \decodedPacket[5][38] ,
         \decodedPacket[5][37] , \decodedPacket[5][4] , \decodedPacket[5][3] ,
         \decodedPacket[5][2] , \decodedPacket[5][1] , \decodedPacket[5][0] ,
         \decodedPacket[4][121] , \decodedPacket[4][120] ,
         \decodedPacket[4][119] , \decodedPacket[4][118] ,
         \decodedPacket[4][117] , \decodedPacket[4][116] ,
         \decodedPacket[4][115] , \decodedPacket[4][114] ,
         \decodedPacket[4][113] , \decodedPacket[4][112] ,
         \decodedPacket[4][111] , \decodedPacket[4][110] ,
         \decodedPacket[4][109] , \decodedPacket[4][108] ,
         \decodedPacket[4][107] , \decodedPacket[4][106] ,
         \decodedPacket[4][105] , \decodedPacket[4][104] ,
         \decodedPacket[4][103] , \decodedPacket[4][102] ,
         \decodedPacket[4][101] , \decodedPacket[4][100] ,
         \decodedPacket[4][99] , \decodedPacket[4][98] ,
         \decodedPacket[4][97] , \decodedPacket[4][96] ,
         \decodedPacket[4][95] , \decodedPacket[4][94] ,
         \decodedPacket[4][93] , \decodedPacket[4][92] ,
         \decodedPacket[4][91] , \decodedPacket[4][90] ,
         \decodedPacket[4][89] , \decodedPacket[4][88] ,
         \decodedPacket[4][87] , \decodedPacket[4][86] ,
         \decodedPacket[4][85] , \decodedPacket[4][84] ,
         \decodedPacket[4][83] , \decodedPacket[4][82] ,
         \decodedPacket[4][81] , \decodedPacket[4][80] ,
         \decodedPacket[4][79] , \decodedPacket[4][78] ,
         \decodedPacket[4][77] , \decodedPacket[4][76] ,
         \decodedPacket[4][75] , \decodedPacket[4][74] ,
         \decodedPacket[4][73] , \decodedPacket[4][72] ,
         \decodedPacket[4][71] , \decodedPacket[4][70] ,
         \decodedPacket[4][69] , \decodedPacket[4][68] ,
         \decodedPacket[4][67] , \decodedPacket[4][66] ,
         \decodedPacket[4][65] , \decodedPacket[4][64] ,
         \decodedPacket[4][63] , \decodedPacket[4][62] ,
         \decodedPacket[4][61] , \decodedPacket[4][60] ,
         \decodedPacket[4][59] , \decodedPacket[4][58] ,
         \decodedPacket[4][57] , \decodedPacket[4][56] ,
         \decodedPacket[4][55] , \decodedPacket[4][54] ,
         \decodedPacket[4][53] , \decodedPacket[4][52] ,
         \decodedPacket[4][51] , \decodedPacket[4][50] ,
         \decodedPacket[4][49] , \decodedPacket[4][48] ,
         \decodedPacket[4][47] , \decodedPacket[4][46] ,
         \decodedPacket[4][45] , \decodedPacket[4][44] ,
         \decodedPacket[4][43] , \decodedPacket[4][42] ,
         \decodedPacket[4][41] , \decodedPacket[4][40] ,
         \decodedPacket[4][39] , \decodedPacket[4][38] ,
         \decodedPacket[4][37] , \decodedPacket[4][36] ,
         \decodedPacket[4][35] , \decodedPacket[4][34] ,
         \decodedPacket[4][33] , \decodedPacket[4][32] ,
         \decodedPacket[4][31] , \decodedPacket[4][30] ,
         \decodedPacket[4][29] , \decodedPacket[4][28] ,
         \decodedPacket[4][27] , \decodedPacket[4][26] ,
         \decodedPacket[4][25] , \decodedPacket[4][24] ,
         \decodedPacket[4][23] , \decodedPacket[4][22] ,
         \decodedPacket[4][21] , \decodedPacket[4][20] ,
         \decodedPacket[4][19] , \decodedPacket[4][18] ,
         \decodedPacket[4][17] , \decodedPacket[4][16] ,
         \decodedPacket[4][15] , \decodedPacket[4][14] ,
         \decodedPacket[4][13] , \decodedPacket[4][12] ,
         \decodedPacket[4][11] , \decodedPacket[4][10] , \decodedPacket[4][9] ,
         \decodedPacket[4][8] , \decodedPacket[4][7] , \decodedPacket[4][6] ,
         \decodedPacket[4][5] , \decodedPacket[4][4] , \decodedPacket[4][3] ,
         \decodedPacket[4][2] , \decodedPacket[4][1] , \decodedPacket[4][0] ,
         \decodedPacket[3][120] , \decodedPacket[3][119] ,
         \decodedPacket[3][118] , \decodedPacket[3][116] ,
         \decodedPacket[3][115] , \decodedPacket[3][114] ,
         \decodedPacket[3][113] , \decodedPacket[3][112] ,
         \decodedPacket[3][111] , \decodedPacket[3][110] ,
         \decodedPacket[3][109] , \decodedPacket[3][108] ,
         \decodedPacket[3][107] , \decodedPacket[3][106] ,
         \decodedPacket[3][105] , \decodedPacket[3][104] ,
         \decodedPacket[3][103] , \decodedPacket[3][102] ,
         \decodedPacket[3][101] , \decodedPacket[3][100] ,
         \decodedPacket[3][99] , \decodedPacket[3][98] ,
         \decodedPacket[3][97] , \decodedPacket[3][96] ,
         \decodedPacket[3][95] , \decodedPacket[3][94] ,
         \decodedPacket[3][93] , \decodedPacket[3][92] ,
         \decodedPacket[3][91] , \decodedPacket[3][90] ,
         \decodedPacket[3][89] , \decodedPacket[3][88] ,
         \decodedPacket[3][87] , \decodedPacket[3][86] ,
         \decodedPacket[3][85] , \decodedPacket[3][84] ,
         \decodedPacket[3][83] , \decodedPacket[3][82] ,
         \decodedPacket[3][81] , \decodedPacket[3][80] ,
         \decodedPacket[3][79] , \decodedPacket[3][78] ,
         \decodedPacket[3][77] , \decodedPacket[3][76] ,
         \decodedPacket[3][75] , \decodedPacket[3][74] ,
         \decodedPacket[3][73] , \decodedPacket[3][72] ,
         \decodedPacket[3][71] , \decodedPacket[3][70] ,
         \decodedPacket[3][69] , \decodedPacket[3][68] ,
         \decodedPacket[3][67] , \decodedPacket[3][66] ,
         \decodedPacket[3][65] , \decodedPacket[3][64] ,
         \decodedPacket[3][63] , \decodedPacket[3][62] ,
         \decodedPacket[3][61] , \decodedPacket[3][60] ,
         \decodedPacket[3][59] , \decodedPacket[3][58] ,
         \decodedPacket[3][57] , \decodedPacket[3][56] ,
         \decodedPacket[3][55] , \decodedPacket[3][54] ,
         \decodedPacket[3][53] , \decodedPacket[3][52] ,
         \decodedPacket[3][51] , \decodedPacket[3][50] ,
         \decodedPacket[3][49] , \decodedPacket[3][48] ,
         \decodedPacket[3][47] , \decodedPacket[3][46] ,
         \decodedPacket[3][45] , \decodedPacket[3][44] ,
         \decodedPacket[3][43] , \decodedPacket[3][42] ,
         \decodedPacket[3][41] , \decodedPacket[3][40] ,
         \decodedPacket[3][39] , \decodedPacket[3][38] ,
         \decodedPacket[3][37] , \decodedPacket[3][4] , \decodedPacket[3][3] ,
         \decodedPacket[3][2] , \decodedPacket[3][1] , \decodedPacket[3][0] ,
         \decodedPacket[2][121] , \decodedPacket[2][120] ,
         \decodedPacket[2][119] , \decodedPacket[2][118] ,
         \decodedPacket[2][117] , \decodedPacket[2][116] ,
         \decodedPacket[2][115] , \decodedPacket[2][114] ,
         \decodedPacket[2][113] , \decodedPacket[2][112] ,
         \decodedPacket[2][111] , \decodedPacket[2][110] ,
         \decodedPacket[2][109] , \decodedPacket[2][108] ,
         \decodedPacket[2][107] , \decodedPacket[2][106] ,
         \decodedPacket[2][105] , \decodedPacket[2][104] ,
         \decodedPacket[2][103] , \decodedPacket[2][102] ,
         \decodedPacket[2][101] , \decodedPacket[2][100] ,
         \decodedPacket[2][99] , \decodedPacket[2][98] ,
         \decodedPacket[2][97] , \decodedPacket[2][96] ,
         \decodedPacket[2][95] , \decodedPacket[2][94] ,
         \decodedPacket[2][93] , \decodedPacket[2][92] ,
         \decodedPacket[2][91] , \decodedPacket[2][90] ,
         \decodedPacket[2][89] , \decodedPacket[2][88] ,
         \decodedPacket[2][87] , \decodedPacket[2][86] ,
         \decodedPacket[2][85] , \decodedPacket[2][84] ,
         \decodedPacket[2][83] , \decodedPacket[2][82] ,
         \decodedPacket[2][81] , \decodedPacket[2][80] ,
         \decodedPacket[2][79] , \decodedPacket[2][78] ,
         \decodedPacket[2][77] , \decodedPacket[2][76] ,
         \decodedPacket[2][75] , \decodedPacket[2][74] ,
         \decodedPacket[2][73] , \decodedPacket[2][72] ,
         \decodedPacket[2][71] , \decodedPacket[2][70] ,
         \decodedPacket[2][69] , \decodedPacket[2][68] ,
         \decodedPacket[2][67] , \decodedPacket[2][66] ,
         \decodedPacket[2][65] , \decodedPacket[2][64] ,
         \decodedPacket[2][63] , \decodedPacket[2][62] ,
         \decodedPacket[2][61] , \decodedPacket[2][60] ,
         \decodedPacket[2][59] , \decodedPacket[2][58] ,
         \decodedPacket[2][57] , \decodedPacket[2][56] ,
         \decodedPacket[2][55] , \decodedPacket[2][54] ,
         \decodedPacket[2][53] , \decodedPacket[2][52] ,
         \decodedPacket[2][51] , \decodedPacket[2][50] ,
         \decodedPacket[2][49] , \decodedPacket[2][48] ,
         \decodedPacket[2][47] , \decodedPacket[2][46] ,
         \decodedPacket[2][45] , \decodedPacket[2][44] ,
         \decodedPacket[2][43] , \decodedPacket[2][42] ,
         \decodedPacket[2][41] , \decodedPacket[2][40] ,
         \decodedPacket[2][39] , \decodedPacket[2][38] ,
         \decodedPacket[2][37] , \decodedPacket[2][36] ,
         \decodedPacket[2][35] , \decodedPacket[2][34] ,
         \decodedPacket[2][33] , \decodedPacket[2][32] ,
         \decodedPacket[2][31] , \decodedPacket[2][30] ,
         \decodedPacket[2][29] , \decodedPacket[2][28] ,
         \decodedPacket[2][27] , \decodedPacket[2][26] ,
         \decodedPacket[2][25] , \decodedPacket[2][24] ,
         \decodedPacket[2][23] , \decodedPacket[2][22] ,
         \decodedPacket[2][21] , \decodedPacket[2][20] ,
         \decodedPacket[2][19] , \decodedPacket[2][18] ,
         \decodedPacket[2][17] , \decodedPacket[2][16] ,
         \decodedPacket[2][15] , \decodedPacket[2][14] ,
         \decodedPacket[2][13] , \decodedPacket[2][12] ,
         \decodedPacket[2][11] , \decodedPacket[2][10] , \decodedPacket[2][9] ,
         \decodedPacket[2][8] , \decodedPacket[2][7] , \decodedPacket[2][6] ,
         \decodedPacket[2][5] , \decodedPacket[2][4] , \decodedPacket[2][3] ,
         \decodedPacket[2][2] , \decodedPacket[2][1] , \decodedPacket[2][0] ,
         \decodedPacket[1][120] , \decodedPacket[1][119] ,
         \decodedPacket[1][118] , \decodedPacket[1][116] ,
         \decodedPacket[1][115] , \decodedPacket[1][114] ,
         \decodedPacket[1][113] , \decodedPacket[1][112] ,
         \decodedPacket[1][111] , \decodedPacket[1][110] ,
         \decodedPacket[1][109] , \decodedPacket[1][108] ,
         \decodedPacket[1][107] , \decodedPacket[1][106] ,
         \decodedPacket[1][105] , \decodedPacket[1][104] ,
         \decodedPacket[1][103] , \decodedPacket[1][102] ,
         \decodedPacket[1][101] , \decodedPacket[1][100] ,
         \decodedPacket[1][99] , \decodedPacket[1][98] ,
         \decodedPacket[1][97] , \decodedPacket[1][96] ,
         \decodedPacket[1][95] , \decodedPacket[1][94] ,
         \decodedPacket[1][93] , \decodedPacket[1][92] ,
         \decodedPacket[1][91] , \decodedPacket[1][90] ,
         \decodedPacket[1][89] , \decodedPacket[1][88] ,
         \decodedPacket[1][87] , \decodedPacket[1][86] ,
         \decodedPacket[1][85] , \decodedPacket[1][84] ,
         \decodedPacket[1][83] , \decodedPacket[1][82] ,
         \decodedPacket[1][81] , \decodedPacket[1][80] ,
         \decodedPacket[1][79] , \decodedPacket[1][78] ,
         \decodedPacket[1][77] , \decodedPacket[1][76] ,
         \decodedPacket[1][75] , \decodedPacket[1][74] ,
         \decodedPacket[1][73] , \decodedPacket[1][72] ,
         \decodedPacket[1][71] , \decodedPacket[1][70] ,
         \decodedPacket[1][69] , \decodedPacket[1][68] ,
         \decodedPacket[1][67] , \decodedPacket[1][66] ,
         \decodedPacket[1][65] , \decodedPacket[1][64] ,
         \decodedPacket[1][63] , \decodedPacket[1][62] ,
         \decodedPacket[1][61] , \decodedPacket[1][60] ,
         \decodedPacket[1][59] , \decodedPacket[1][58] ,
         \decodedPacket[1][57] , \decodedPacket[1][56] ,
         \decodedPacket[1][55] , \decodedPacket[1][54] ,
         \decodedPacket[1][53] , \decodedPacket[1][52] ,
         \decodedPacket[1][51] , \decodedPacket[1][50] ,
         \decodedPacket[1][49] , \decodedPacket[1][48] ,
         \decodedPacket[1][47] , \decodedPacket[1][46] ,
         \decodedPacket[1][45] , \decodedPacket[1][44] ,
         \decodedPacket[1][43] , \decodedPacket[1][42] ,
         \decodedPacket[1][41] , \decodedPacket[1][40] ,
         \decodedPacket[1][39] , \decodedPacket[1][38] ,
         \decodedPacket[1][37] , \decodedPacket[1][4] , \decodedPacket[1][3] ,
         \decodedPacket[1][2] , \decodedPacket[1][1] , \decodedPacket[1][0] ,
         \decodedPacket[0][121] , \decodedPacket[0][120] ,
         \decodedPacket[0][119] , \decodedPacket[0][118] ,
         \decodedPacket[0][117] , \decodedPacket[0][116] ,
         \decodedPacket[0][115] , \decodedPacket[0][114] ,
         \decodedPacket[0][113] , \decodedPacket[0][112] ,
         \decodedPacket[0][111] , \decodedPacket[0][110] ,
         \decodedPacket[0][109] , \decodedPacket[0][108] ,
         \decodedPacket[0][107] , \decodedPacket[0][106] ,
         \decodedPacket[0][105] , \decodedPacket[0][104] ,
         \decodedPacket[0][103] , \decodedPacket[0][102] ,
         \decodedPacket[0][101] , \decodedPacket[0][100] ,
         \decodedPacket[0][99] , \decodedPacket[0][98] ,
         \decodedPacket[0][97] , \decodedPacket[0][96] ,
         \decodedPacket[0][95] , \decodedPacket[0][94] ,
         \decodedPacket[0][93] , \decodedPacket[0][92] ,
         \decodedPacket[0][91] , \decodedPacket[0][90] ,
         \decodedPacket[0][89] , \decodedPacket[0][88] ,
         \decodedPacket[0][87] , \decodedPacket[0][86] ,
         \decodedPacket[0][85] , \decodedPacket[0][84] ,
         \decodedPacket[0][83] , \decodedPacket[0][82] ,
         \decodedPacket[0][81] , \decodedPacket[0][80] ,
         \decodedPacket[0][79] , \decodedPacket[0][78] ,
         \decodedPacket[0][77] , \decodedPacket[0][76] ,
         \decodedPacket[0][75] , \decodedPacket[0][74] ,
         \decodedPacket[0][73] , \decodedPacket[0][72] ,
         \decodedPacket[0][71] , \decodedPacket[0][70] ,
         \decodedPacket[0][69] , \decodedPacket[0][68] ,
         \decodedPacket[0][67] , \decodedPacket[0][66] ,
         \decodedPacket[0][65] , \decodedPacket[0][64] ,
         \decodedPacket[0][63] , \decodedPacket[0][62] ,
         \decodedPacket[0][61] , \decodedPacket[0][60] ,
         \decodedPacket[0][59] , \decodedPacket[0][58] ,
         \decodedPacket[0][57] , \decodedPacket[0][56] ,
         \decodedPacket[0][55] , \decodedPacket[0][54] ,
         \decodedPacket[0][53] , \decodedPacket[0][52] ,
         \decodedPacket[0][51] , \decodedPacket[0][50] ,
         \decodedPacket[0][49] , \decodedPacket[0][48] ,
         \decodedPacket[0][47] , \decodedPacket[0][46] ,
         \decodedPacket[0][45] , \decodedPacket[0][44] ,
         \decodedPacket[0][43] , \decodedPacket[0][42] ,
         \decodedPacket[0][41] , \decodedPacket[0][40] ,
         \decodedPacket[0][39] , \decodedPacket[0][38] ,
         \decodedPacket[0][37] , \decodedPacket[0][36] ,
         \decodedPacket[0][35] , \decodedPacket[0][34] ,
         \decodedPacket[0][33] , \decodedPacket[0][32] ,
         \decodedPacket[0][31] , \decodedPacket[0][30] ,
         \decodedPacket[0][29] , \decodedPacket[0][28] ,
         \decodedPacket[0][27] , \decodedPacket[0][26] ,
         \decodedPacket[0][25] , \decodedPacket[0][24] ,
         \decodedPacket[0][23] , \decodedPacket[0][22] ,
         \decodedPacket[0][21] , \decodedPacket[0][20] ,
         \decodedPacket[0][19] , \decodedPacket[0][18] ,
         \decodedPacket[0][17] , \decodedPacket[0][16] ,
         \decodedPacket[0][15] , \decodedPacket[0][14] ,
         \decodedPacket[0][13] , \decodedPacket[0][12] ,
         \decodedPacket[0][11] , \decodedPacket[0][10] , \decodedPacket[0][9] ,
         \decodedPacket[0][8] , \decodedPacket[0][7] , \decodedPacket[0][6] ,
         \decodedPacket[0][5] , \decodedPacket[0][4] , \decodedPacket[0][3] ,
         \decodedPacket[0][2] , \decodedPacket[0][1] , \decodedPacket[0][0] ,
         N389, N1068, N1069, N1070, N2172, N2173, N2174, N2175, N4308, N4309,
         N4310, N4311, N4312, N6444, N6445, N6446, N6447, N6448, N6449, N8580,
         N8581, N8582, N8583, N8584, N8585, N9669, N9670, N9671, N9672, N9673,
         N9674, N9675, N9676, N9677, N9678, N9679, N9680, N9681, N9682, N9683,
         N9684, N9685, N9686, N9687, N9688, N9689, N9690, N9691, N9692, N9693,
         N9694, N9695, N9696, N9697, N9698, N9699, N9700, N9701, N9702, N9703,
         N9704, N9705, N9706, N9707, N9708, N9709, N9710, N9711, N9712, N9713,
         N9714, N9715, N9716, N9718, N9719, N9720, N9721, N9722, N9723, N9724,
         N9725, N9726, N9727, N9728, N9729, N9730, N9731, N9732, N9733, N9734,
         N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9743, N9744,
         N9745, N9746, N9747, N9748, N9749, N9750, N9751, N9752, N9753, N9754,
         N9755, N9756, N9757, N9758, N9759, N9760, N9761, N9762, N9763, N9764,
         N9765, N9766, N9768, N9769, N9770, N9771, N9772, N9773, N9774, N9775,
         N9776, N9777, N9778, N9779, N9780, N9781, N9782, N9783, N9784, N9785,
         N9786, N9787, N9788, N9789, N9790, N9791, N9792, N9798, N9799, N9800,
         N9801, N9802, N9803, N9804, N9805, N9806, N9807, N9808, N9809, N9810,
         N9811, N9812, N9813, N9814, N9815, N9816, N9817, N9818, N9819, N9820,
         N9821, N9822, N9823, N9824, N9825, N9826, N9827, N9828, N9829, N9830,
         N9831, N9832, N9833, N9834, N9835, N9836, N9837, N9838, N9839, N9840,
         N9841, N9842, N9843, N9844, N9845, N9846, N9848, N9849, N9850, N9851,
         N9852, N9853, N9854, N9855, N9856, N9857, N9858, N9859, N9860, N9861,
         N9862, N9863, N9864, N9865, N9866, N9867, N9868, N9869, N9870, N9871,
         N9872, N9873, N9874, N9875, N9876, N9877, N9878, N9879, N9880, N9881,
         N9882, N9883, N9884, N9885, N9886, N9887, N9888, N9889, N9890, N9891,
         N9892, N9893, N9894, N9895, N9896, N9898, N9900, N9901, N9902, N9903,
         N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9912, N9913,
         N9914, N9915, N9916, N9917, N9918, N9919, N9920, N9921, N9922, N9928,
         N9929, N9930, N9931, N9932, N9933, N9934, N9935, N9936, N9937, N9938,
         N9939, N9940, N9941, N9942, N9943, N9944, N9945, N9946, N9947, N9948,
         N9949, N9950, N9951, N9952, N9953, N9954, N9955, N9956, N9957, N9958,
         N9959, N9960, N9961, N9962, N9963, N9964, N9965, N9966, N9967, N9968,
         N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9978, N9979,
         N9980, N9981, N9982, N9983, N9984, N9985, N9986, N9987, N9988, N9989,
         N9990, N9991, N9992, N9993, N9994, N9995, N9996, N9997, N9998, N9999,
         N10000, N10001, N10002, N10003, N10004, N10005, N10006, N10007,
         N10008, N10009, N10010, N10011, N10012, N10013, N10014, N10015,
         N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023,
         N10024, N10025, N10026, N10028, N10030, N10031, N10032, N10033,
         N10034, N10035, N10036, N10037, N10038, N10039, N10040, N10041,
         N10042, N10043, N10044, N10045, N10046, N10047, N10048, N10049,
         N10050, N10051, N10052, N10058, N10059, N10060, N10061, N10062,
         N10063, N10064, N10065, N10066, N10067, N10068, N10069, N10070,
         N10071, N10072, N10073, N10074, N10075, N10076, N10077, N10078,
         N10079, N10080, N10081, N10082, N10083, N10084, N10085, N10086,
         N10087, N10088, N10089, N10090, N10091, N10092, N10093, N10094,
         N10095, N10096, N10097, N10098, N10099, N10100, N10101, N10102,
         N10103, N10104, N10105, N10106, N10108, N10109, N10110, N10111,
         N10112, N10113, N10114, N10115, N10116, N10117, N10118, N10119,
         N10120, N10121, N10122, N10123, N10124, N10125, N10126, N10127,
         N10128, N10129, N10130, N10131, N10132, N10133, N10134, N10135,
         N10136, N10137, N10138, N10139, N10140, N10141, N10142, N10143,
         N10144, N10145, N10146, N10147, N10148, N10149, N10150, N10151,
         N10152, N10153, N10154, N10155, N10156, N10158, N10160, N10161,
         N10162, N10163, N10164, N10165, N10166, N10167, N10168, N10169,
         N10170, N10171, N10172, N10173, N10174, N10175, N10176, N10177,
         N10178, N10179, N10180, N10181, N10182, N10188, N10189, N10190,
         N10191, N10192, N10193, N10194, N10195, N10196, N10197, N10198,
         N10199, N10200, N10201, N10202, N10203, N10204, N10205, N10206,
         N10207, N10208, N10209, N10210, N10211, N10212, N10213, N10214,
         N10215, N10216, N10217, N10218, N10219, N10220, N10221, N10222,
         N10223, N10224, N10225, N10226, N10227, N10228, N10229, N10230,
         N10231, N10232, N10233, N10234, N10235, N10236, N10238, N10239,
         N10240, N10241, N10242, N10243, N10244, N10245, N10246, N10247,
         N10248, N10249, N10250, N10251, N10252, N10253, N10254, N10255,
         N10256, N10257, N10258, N10259, N10260, N10261, N10262, N10263,
         N10264, N10265, N10266, N10267, N10268, N10269, N10270, N10271,
         N10272, N10273, N10274, N10275, N10276, N10277, N10278, N10279,
         N10280, N10281, N10282, N10283, N10284, N10285, N10286, N10288,
         N10290, N10291, N10292, N10293, N10294, N10295, N10296, N10297,
         N10298, N10299, N10300, N10301, N10302, N10303, N10304, N10305,
         N10306, N10307, N10308, N10309, N10310, N10311, N10312, N10318,
         N10319, N10320, N10321, N10322, N10323, N10324, N10325, N10326,
         N10327, N10328, N10329, N10330, N10331, N10332, N10333, N10334,
         N10335, N10336, N10337, N10338, N10339, N10340, N10341, N10342,
         N10343, N10344, N10345, N10346, N10347, N10348, N10349, N10350,
         N10351, N10352, N10353, N10354, N10355, N10356, N10357, N10358,
         N10359, N10360, N10361, N10362, N10363, N10364, N10365, N10366,
         N10368, N10369, N10370, N10371, N10372, N10373, N10374, N10375,
         N10376, N10377, N10378, N10379, N10380, N10381, N10382, N10383,
         N10384, N10385, N10386, N10387, N10388, N10389, N10390, N10391,
         N10392, N10393, N10394, N10395, N10396, N10397, N10398, N10399,
         N10400, N10401, N10402, N10403, N10404, N10405, N10406, N10407,
         N10408, N10409, N10410, N10411, N10412, N10413, N10414, N10415,
         N10416, N10418, N10420, N10421, N10422, N10423, N10424, N10425,
         N10426, N10427, N10428, N10429, N10430, N10431, N10432, N10433,
         N10434, N10435, N10436, N10437, N10438, N10439, N10440, N10441,
         N10442, N10448, N10449, N10450, N10451, N10452, N10453, N10454,
         N10455, N10456, N10457, N10458, N10459, N10460, N10461, N10462,
         N10463, N10464, N10465, N10466, N10467, N10468, N10469, N10470,
         N10471, N10472, N10473, N10474, N10475, N10476, N10477, N10478,
         N10479, N10480, N10481, N10482, N10483, N10484, N10485, N10486,
         N10487, N10488, N10489, N10490, N10491, N10492, N10493, N10494,
         N10495, N10496, N10498, N10499, N10500, N10501, N10502, N10503,
         N10504, N10505, N10506, N10507, N10508, N10509, N10510, N10511,
         N10512, N10513, N10514, N10515, N10516, N10517, N10518, N10519,
         N10520, N10521, N10522, N10523, N10524, N10525, N10526, N10527,
         N10528, N10529, N10530, N10531, N10532, N10533, N10534, N10535,
         N10536, N10537, N10538, N10539, N10540, N10541, N10542, N10543,
         N10544, N10545, N10546, N10548, N10550, N10551, N10552, N10553,
         N10554, N10555, N10556, N10557, N10558, N10559, N10560, N10561,
         N10562, N10563, N10564, N10565, N10566, N10567, N10568, N10569,
         N10570, N10571, N10572, N10578, N10579, N10580, N10581, N10582,
         N10583, N10584, N10585, N10586, N10587, N10588, N10589, N10590,
         N10591, N10592, N10593, N10594, N10595, N10596, N10597, N10598,
         N10599, N10600, N10601, N10602, N10603, N10604, N10605, N10606,
         N10607, N10608, N10609, N10610, N10611, N10612, N10613, N10614,
         N10615, N10616, N10617, N10618, N10619, N10620, N10621, N10622,
         N10623, N10624, N10625, N10626, N10628, N10629, N10630, N10631,
         N10632, N10633, N10634, N10635, N10636, N10637, N10638, N10639,
         N10640, N10641, N10642, N10643, N10644, N10645, N10646, N10647,
         N10648, N10649, N10650, N10651, N10652, N10653, N10654, N10655,
         N10656, N10657, N10658, N10659, N10660, N10661, N10662, N10663,
         N10664, N10665, N10666, N10667, N10668, N10669, N10670, N10671,
         N10672, N10673, N10674, N10675, N10676, N10678, N10680, N10681,
         N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689,
         N10690, N10691, N10692, N10693, N10694, N10695, N10696, N10697,
         N10698, N10699, N10700, N10701, N10702, n825, n826, n827, n828, n830,
         n831, n832, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n969, n970, n971, n973, n974, n975, n977,
         n978, n979, n981, n982, n983, n985, n986, n987, n989, n990, n991,
         n993, n994, n995, n997, n998, n999, n1001, n1002, n1003, n1005, n1006,
         n1007, n1009, n1010, n1011, n1013, n1014, n1015, n1017, n1018, n1019,
         n1021, n1022, n1023, n1025, n1026, n1027, n1029, n1030, n1031, n1033,
         n1034, n1035, n1037, n1038, n1039, n1041, n1042, n1043, n1045, n1046,
         n1047, n1049, n1050, n1051, n1053, n1054, n1055, n1057, n1058, n1059,
         n1061, n1062, n1063, n1065, n1066, n1067, n1069, n1070, n1071, n1073,
         n1074, n1075, n1077, n1078, n1079, n1081, n1082, n1083, n1085, n1086,
         n1087, n1089, n1090, n1091, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1116, n1124, n1140, n1141,
         n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1163, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1568, n1570, n1571, n1573, n1575, n1576, n1578, n1580, n1581,
         n1583, n1585, n1586, n1588, n1590, n1591, n1593, n1595, n1596, n1598,
         n1600, n1601, n1603, n1605, n1606, n1608, n1610, n1611, n1613, n1615,
         n1616, n1618, n1620, n1621, n1623, n1625, n1626, n1628, n1630, n1631,
         n1633, n1635, n1636, n1638, n1640, n1641, n1643, n1645, n1646, n1648,
         n1650, n1651, n1653, n1655, n1656, n1658, n1660, n1661, n1663, n1665,
         n1666, n1668, n1670, n1671, n1673, n1675, n1676, n1678, n1680, n1681,
         n1683, n1685, n1686, n1688, n1690, n1691, n1693, n1695, n1696, n1698,
         n1700, n1701, n1703, n1705, n1706, n1708, n1710, n1711, n1713, n1715,
         n1716, n1718, n1720, n1721, n1723, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1752, n1753, n1754, n1755, n1757, n1759, n1763, n1767, n1768,
         n1787, n1788, n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1814, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2300, n2302,
         n2303, n2304, n2306, n2308, n2309, n2310, n2312, n2314, n2315, n2316,
         n2318, n2320, n2321, n2322, n2324, n2326, n2327, n2328, n2330, n2332,
         n2333, n2334, n2336, n2338, n2339, n2340, n2342, n2344, n2345, n2346,
         n2348, n2350, n2351, n2352, n2354, n2356, n2357, n2358, n2360, n2362,
         n2363, n2364, n2366, n2368, n2369, n2370, n2372, n2374, n2375, n2376,
         n2378, n2380, n2381, n2382, n2384, n2386, n2387, n2388, n2390, n2392,
         n2393, n2394, n2396, n2398, n2399, n2400, n2402, n2404, n2405, n2406,
         n2408, n2410, n2411, n2412, n2414, n2416, n2417, n2418, n2420, n2422,
         n2423, n2424, n2426, n2428, n2429, n2430, n2432, n2434, n2435, n2436,
         n2438, n2440, n2441, n2442, n2444, n2446, n2447, n2448, n2450, n2452,
         n2453, n2454, n2456, n2458, n2459, n2460, n2462, n2464, n2465, n2466,
         n2468, n2470, n2471, n2472, n2474, n2476, n2477, n2478, n2480, n2482,
         n2483, n2484, n2486, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2525,
         n2529, n2539, n2540, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2797, n2798, n2800, n2801,
         n2803, n2804, n2806, n2807, n2809, n2810, n2812, n2813, n2815, n2816,
         n2818, n2819, n2821, n2822, n2824, n2825, n2827, n2828, n2830, n2831,
         n2833, n2834, n2836, n2837, n2839, n2840, n2842, n2843, n2845, n2846,
         n2848, n2849, n2851, n2852, n2854, n2855, n2857, n2858, n2860, n2861,
         n2863, n2864, n2866, n2867, n2869, n2870, n2872, n2873, n2875, n2876,
         n2878, n2879, n2881, n2882, n2884, n2885, n2887, n2888, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2912,
         n2914, n2918, n2928, n2929, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3186, n3187, n3189,
         n3190, n3192, n3193, n3195, n3196, n3198, n3199, n3201, n3202, n3204,
         n3205, n3207, n3208, n3210, n3211, n3213, n3214, n3216, n3217, n3219,
         n3220, n3222, n3223, n3225, n3226, n3228, n3229, n3231, n3232, n3234,
         n3235, n3237, n3238, n3240, n3241, n3243, n3244, n3246, n3247, n3249,
         n3250, n3252, n3253, n3255, n3256, n3258, n3259, n3261, n3262, n3264,
         n3265, n3267, n3268, n3270, n3271, n3273, n3274, n3276, n3277, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, n3302, n3312,
         n3313, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3570, n3571, n3573, n3574, n3576, n3577,
         n3579, n3580, n3582, n3583, n3585, n3586, n3588, n3589, n3591, n3592,
         n3594, n3595, n3597, n3598, n3600, n3601, n3603, n3604, n3606, n3607,
         n3609, n3610, n3612, n3613, n3615, n3616, n3618, n3619, n3621, n3622,
         n3624, n3625, n3627, n3628, n3630, n3631, n3633, n3634, n3636, n3637,
         n3639, n3640, n3642, n3643, n3645, n3646, n3648, n3649, n3651, n3652,
         n3654, n3655, n3657, n3658, n3660, n3661, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3682, n3686, n3696, n3697, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3954, n3955, n3957, n3958, n3960, n3961, n3963, n3964, n3966,
         n3967, n3969, n3970, n3972, n3973, n3975, n3976, n3978, n3979, n3981,
         n3982, n3984, n3985, n3987, n3988, n3990, n3991, n3993, n3994, n3996,
         n3997, n3999, n4000, n4002, n4003, n4005, n4006, n4008, n4009, n4011,
         n4012, n4014, n4015, n4017, n4018, n4020, n4021, n4023, n4024, n4026,
         n4027, n4029, n4030, n4032, n4033, n4035, n4036, n4038, n4039, n4041,
         n4042, n4044, n4045, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4066, n4070, n4072, n4076, n4090, n4091, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4433, n4434, n4435, n4437, n4438, n4439,
         n4441, n4442, n4443, n4445, n4446, n4447, n4449, n4450, n4451, n4453,
         n4454, n4455, n4457, n4458, n4459, n4461, n4462, n4463, n4465, n4466,
         n4467, n4469, n4470, n4471, n4473, n4474, n4475, n4477, n4478, n4479,
         n4481, n4482, n4483, n4485, n4486, n4487, n4489, n4490, n4491, n4493,
         n4494, n4495, n4497, n4498, n4499, n4501, n4502, n4503, n4505, n4506,
         n4507, n4509, n4510, n4511, n4513, n4514, n4515, n4517, n4518, n4519,
         n4521, n4522, n4523, n4525, n4526, n4527, n4529, n4530, n4531, n4533,
         n4534, n4535, n4537, n4538, n4539, n4541, n4542, n4543, n4545, n4546,
         n4547, n4549, n4550, n4551, n4553, n4554, n4555, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4595,
         n4596, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4837, \add_177_I7_aco/carry[1] ,
         \add_177_I7_aco/carry[2] , \add_177_I7_aco/carry[3] ,
         \add_177_I7_aco/carry[4] , \add_177_I7_aco/carry[5] ,
         \add_177_I6_aco/carry[1] , \add_177_I6_aco/carry[2] ,
         \add_177_I6_aco/carry[3] , \add_177_I6_aco/carry[4] ,
         \add_177_I5_aco/carry[1] , \add_177_I5_aco/carry[2] ,
         \add_177_I5_aco/carry[3] , \add_177_I4_aco/carry[1] ,
         \add_177_I4_aco/carry[2] , \add_177_I3_aco/carry[1] ,
         \add_177_I3_aco/A[0] , \add_177_I3_aco/A[1] , n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459;
  wire   [7:0] decodedPacketValid;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167;

  LATCHX1 \decodedPacket_f_reg[7][121]  ( .CLK(n5931), .D(N10702), .Q(
        decodedPacket7_o[121]) );
  LATCHX1 \decodedPacket_f_reg[7][120]  ( .CLK(n5932), .D(N10701), .Q(
        decodedPacket7_o[120]) );
  LATCHX1 \decodedPacket_f_reg[7][119]  ( .CLK(n5936), .D(N10700), .Q(
        decodedPacket7_o[119]) );
  LATCHX1 \decodedPacket_f_reg[7][118]  ( .CLK(n5936), .D(N10699), .Q(
        decodedPacket7_o[118]) );
  LATCHX1 \decodedPacket_f_reg[7][117]  ( .CLK(n5936), .D(N10698), .Q(
        decodedPacket7_o[117]) );
  LATCHX1 \decodedPacket_f_reg[7][116]  ( .CLK(n5936), .D(N10697), .Q(
        decodedPacket7_o[116]) );
  LATCHX1 \decodedPacket_f_reg[7][115]  ( .CLK(n5936), .D(N10696), .Q(
        decodedPacket7_o[115]) );
  LATCHX1 \decodedPacket_f_reg[7][114]  ( .CLK(n5936), .D(N10695), .Q(
        decodedPacket7_o[114]) );
  LATCHX1 \decodedPacket_f_reg[7][113]  ( .CLK(n5936), .D(N10694), .Q(
        decodedPacket7_o[113]) );
  LATCHX1 \decodedPacket_f_reg[7][112]  ( .CLK(n5936), .D(N10693), .Q(
        decodedPacket7_o[112]) );
  LATCHX1 \decodedPacket_f_reg[7][111]  ( .CLK(n5936), .D(N10692), .Q(
        decodedPacket7_o[111]) );
  LATCHX1 \decodedPacket_f_reg[7][110]  ( .CLK(n5936), .D(N10691), .Q(
        decodedPacket7_o[110]) );
  LATCHX1 \decodedPacket_f_reg[7][109]  ( .CLK(n5936), .D(N10690), .Q(
        decodedPacket7_o[109]) );
  LATCHX1 \decodedPacket_f_reg[7][108]  ( .CLK(n5936), .D(N10689), .Q(
        decodedPacket7_o[108]) );
  LATCHX1 \decodedPacket_f_reg[7][107]  ( .CLK(n5935), .D(N10688), .Q(
        decodedPacket7_o[107]) );
  LATCHX1 \decodedPacket_f_reg[7][106]  ( .CLK(n5935), .D(N10687), .Q(
        decodedPacket7_o[106]) );
  LATCHX1 \decodedPacket_f_reg[7][105]  ( .CLK(n5935), .D(N10686), .Q(
        decodedPacket7_o[105]) );
  LATCHX1 \decodedPacket_f_reg[7][104]  ( .CLK(n5935), .D(N10685), .Q(
        decodedPacket7_o[104]) );
  LATCHX1 \decodedPacket_f_reg[7][103]  ( .CLK(n5935), .D(N10684), .Q(
        decodedPacket7_o[103]) );
  LATCHX1 \decodedPacket_f_reg[7][102]  ( .CLK(n5935), .D(N10683), .Q(
        decodedPacket7_o[102]) );
  LATCHX1 \decodedPacket_f_reg[7][101]  ( .CLK(n5935), .D(N10682), .Q(
        decodedPacket7_o[101]) );
  LATCHX1 \decodedPacket_f_reg[7][100]  ( .CLK(n5935), .D(N10681), .Q(
        decodedPacket7_o[100]) );
  LATCHX1 \decodedPacket_f_reg[7][99]  ( .CLK(n5935), .D(N10680), .Q(
        decodedPacket7_o[99]) );
  LATCHX1 \decodedPacket_f_reg[7][98]  ( .CLK(n5935), .D(N10678), .Q(
        decodedPacket7_o[98]) );
  LATCHX1 \decodedPacket_f_reg[7][97]  ( .CLK(n5935), .D(N10676), .Q(
        decodedPacket7_o[97]) );
  LATCHX1 \decodedPacket_f_reg[7][96]  ( .CLK(n5935), .D(N10675), .Q(
        decodedPacket7_o[96]) );
  LATCHX1 \decodedPacket_f_reg[7][95]  ( .CLK(n5934), .D(N10674), .Q(
        decodedPacket7_o[95]) );
  LATCHX1 \decodedPacket_f_reg[7][94]  ( .CLK(n5934), .D(N10673), .Q(
        decodedPacket7_o[94]) );
  LATCHX1 \decodedPacket_f_reg[7][93]  ( .CLK(n5934), .D(N10672), .Q(
        decodedPacket7_o[93]) );
  LATCHX1 \decodedPacket_f_reg[7][92]  ( .CLK(n5934), .D(N10671), .Q(
        decodedPacket7_o[92]) );
  LATCHX1 \decodedPacket_f_reg[7][91]  ( .CLK(n5934), .D(N10670), .Q(
        decodedPacket7_o[91]) );
  LATCHX1 \decodedPacket_f_reg[7][90]  ( .CLK(n5934), .D(N10669), .Q(
        decodedPacket7_o[90]) );
  LATCHX1 \decodedPacket_f_reg[7][89]  ( .CLK(n5934), .D(N10668), .Q(
        decodedPacket7_o[89]) );
  LATCHX1 \decodedPacket_f_reg[7][88]  ( .CLK(n5934), .D(N10667), .Q(
        decodedPacket7_o[88]) );
  LATCHX1 \decodedPacket_f_reg[7][87]  ( .CLK(n5934), .D(N10666), .Q(
        decodedPacket7_o[87]) );
  LATCHX1 \decodedPacket_f_reg[7][86]  ( .CLK(n5934), .D(N10665), .Q(
        decodedPacket7_o[86]) );
  LATCHX1 \decodedPacket_f_reg[7][85]  ( .CLK(n5934), .D(N10664), .Q(
        decodedPacket7_o[85]) );
  LATCHX1 \decodedPacket_f_reg[7][84]  ( .CLK(n5934), .D(N10663), .Q(
        decodedPacket7_o[84]) );
  LATCHX1 \decodedPacket_f_reg[7][83]  ( .CLK(n5933), .D(N10662), .Q(
        decodedPacket7_o[83]) );
  LATCHX1 \decodedPacket_f_reg[7][82]  ( .CLK(n5933), .D(N10661), .Q(
        decodedPacket7_o[82]) );
  LATCHX1 \decodedPacket_f_reg[7][81]  ( .CLK(n5933), .D(N10660), .Q(
        decodedPacket7_o[81]) );
  LATCHX1 \decodedPacket_f_reg[7][80]  ( .CLK(n5933), .D(N10659), .Q(
        decodedPacket7_o[80]) );
  LATCHX1 \decodedPacket_f_reg[7][79]  ( .CLK(n5933), .D(N10658), .Q(
        decodedPacket7_o[79]) );
  LATCHX1 \decodedPacket_f_reg[7][78]  ( .CLK(n5933), .D(N10657), .Q(
        decodedPacket7_o[78]) );
  LATCHX1 \decodedPacket_f_reg[7][77]  ( .CLK(n5933), .D(N10656), .Q(
        decodedPacket7_o[77]) );
  LATCHX1 \decodedPacket_f_reg[7][76]  ( .CLK(n5933), .D(N10655), .Q(
        decodedPacket7_o[76]) );
  LATCHX1 \decodedPacket_f_reg[7][75]  ( .CLK(n5933), .D(N10654), .Q(
        decodedPacket7_o[75]) );
  LATCHX1 \decodedPacket_f_reg[7][74]  ( .CLK(n5933), .D(N10653), .Q(
        decodedPacket7_o[74]) );
  LATCHX1 \decodedPacket_f_reg[7][73]  ( .CLK(n5933), .D(N10652), .Q(
        decodedPacket7_o[73]) );
  LATCHX1 \decodedPacket_f_reg[7][72]  ( .CLK(n5933), .D(N10651), .Q(
        decodedPacket7_o[72]) );
  LATCHX1 \decodedPacket_f_reg[7][71]  ( .CLK(n5932), .D(N10650), .Q(
        decodedPacket7_o[71]) );
  LATCHX1 \decodedPacket_f_reg[7][70]  ( .CLK(n5932), .D(N10649), .Q(
        decodedPacket7_o[70]) );
  LATCHX1 \decodedPacket_f_reg[7][69]  ( .CLK(n5932), .D(N10648), .Q(
        decodedPacket7_o[69]) );
  LATCHX1 \decodedPacket_f_reg[7][68]  ( .CLK(n5932), .D(N10647), .Q(
        decodedPacket7_o[68]) );
  LATCHX1 \decodedPacket_f_reg[7][67]  ( .CLK(n5932), .D(N10646), .Q(
        decodedPacket7_o[67]) );
  LATCHX1 \decodedPacket_f_reg[7][66]  ( .CLK(n5932), .D(N10645), .Q(
        decodedPacket7_o[66]) );
  LATCHX1 \decodedPacket_f_reg[7][65]  ( .CLK(n5932), .D(N10644), .Q(
        decodedPacket7_o[65]) );
  LATCHX1 \decodedPacket_f_reg[7][64]  ( .CLK(n5932), .D(N10643), .Q(
        decodedPacket7_o[64]) );
  LATCHX1 \decodedPacket_f_reg[7][63]  ( .CLK(n5932), .D(N10642), .Q(
        decodedPacket7_o[63]) );
  LATCHX1 \decodedPacket_f_reg[7][62]  ( .CLK(n5932), .D(N10641), .Q(
        decodedPacket7_o[62]) );
  LATCHX1 \decodedPacket_f_reg[7][61]  ( .CLK(n5932), .D(N10640), .Q(
        decodedPacket7_o[61]) );
  LATCHX1 \decodedPacket_f_reg[7][60]  ( .CLK(n5932), .D(N10639), .Q(
        decodedPacket7_o[60]) );
  LATCHX1 \decodedPacket_f_reg[7][59]  ( .CLK(n5931), .D(N10638), .Q(
        decodedPacket7_o[59]) );
  LATCHX1 \decodedPacket_f_reg[7][58]  ( .CLK(n5931), .D(N10637), .Q(
        decodedPacket7_o[58]) );
  LATCHX1 \decodedPacket_f_reg[7][57]  ( .CLK(n5931), .D(N10636), .Q(
        decodedPacket7_o[57]) );
  LATCHX1 \decodedPacket_f_reg[7][56]  ( .CLK(n5931), .D(N10635), .Q(
        decodedPacket7_o[56]) );
  LATCHX1 \decodedPacket_f_reg[7][55]  ( .CLK(n5931), .D(N10634), .Q(
        decodedPacket7_o[55]) );
  LATCHX1 \decodedPacket_f_reg[7][54]  ( .CLK(n5931), .D(N10633), .Q(
        decodedPacket7_o[54]) );
  LATCHX1 \decodedPacket_f_reg[7][53]  ( .CLK(n5931), .D(N10632), .Q(
        decodedPacket7_o[53]) );
  LATCHX1 \decodedPacket_f_reg[7][52]  ( .CLK(n5931), .D(N10631), .Q(
        decodedPacket7_o[52]) );
  LATCHX1 \decodedPacket_f_reg[7][51]  ( .CLK(n5931), .D(N10630), .Q(
        decodedPacket7_o[51]) );
  LATCHX1 \decodedPacket_f_reg[7][50]  ( .CLK(n5931), .D(N10629), .Q(
        decodedPacket7_o[50]) );
  LATCHX1 \decodedPacket_f_reg[7][49]  ( .CLK(n5931), .D(N10628), .Q(
        decodedPacket7_o[49]) );
  LATCHX1 \decodedPacket_f_reg[7][48]  ( .CLK(n5931), .D(N10626), .Q(
        decodedPacket7_o[48]) );
  LATCHX1 \decodedPacket_f_reg[7][47]  ( .CLK(n5930), .D(N10625), .Q(
        decodedPacket7_o[47]) );
  LATCHX1 \decodedPacket_f_reg[7][46]  ( .CLK(n5930), .D(N10624), .Q(
        decodedPacket7_o[46]) );
  LATCHX1 \decodedPacket_f_reg[7][45]  ( .CLK(n5930), .D(N10623), .Q(
        decodedPacket7_o[45]) );
  LATCHX1 \decodedPacket_f_reg[7][44]  ( .CLK(n5930), .D(N10622), .Q(
        decodedPacket7_o[44]) );
  LATCHX1 \decodedPacket_f_reg[7][43]  ( .CLK(n5930), .D(N10621), .Q(
        decodedPacket7_o[43]) );
  LATCHX1 \decodedPacket_f_reg[7][42]  ( .CLK(n5930), .D(N10620), .Q(
        decodedPacket7_o[42]) );
  LATCHX1 \decodedPacket_f_reg[7][41]  ( .CLK(n5930), .D(N10619), .Q(
        decodedPacket7_o[41]) );
  LATCHX1 \decodedPacket_f_reg[7][40]  ( .CLK(n5930), .D(N10618), .Q(
        decodedPacket7_o[40]) );
  LATCHX1 \decodedPacket_f_reg[7][39]  ( .CLK(n5930), .D(N10617), .Q(
        decodedPacket7_o[39]) );
  LATCHX1 \decodedPacket_f_reg[7][38]  ( .CLK(n5930), .D(N10616), .Q(
        decodedPacket7_o[38]) );
  LATCHX1 \decodedPacket_f_reg[7][37]  ( .CLK(n5930), .D(N10615), .Q(
        decodedPacket7_o[37]) );
  LATCHX1 \decodedPacket_f_reg[7][36]  ( .CLK(n5930), .D(N10614), .Q(
        decodedPacket7_o[36]) );
  LATCHX1 \decodedPacket_f_reg[7][35]  ( .CLK(n5929), .D(N10613), .Q(
        decodedPacket7_o[35]) );
  LATCHX1 \decodedPacket_f_reg[7][34]  ( .CLK(n5929), .D(N10612), .Q(
        decodedPacket7_o[34]) );
  LATCHX1 \decodedPacket_f_reg[7][33]  ( .CLK(n5929), .D(N10611), .Q(
        decodedPacket7_o[33]) );
  LATCHX1 \decodedPacket_f_reg[7][32]  ( .CLK(n5929), .D(N10610), .Q(
        decodedPacket7_o[32]) );
  LATCHX1 \decodedPacket_f_reg[7][31]  ( .CLK(n5929), .D(N10609), .Q(
        decodedPacket7_o[31]) );
  LATCHX1 \decodedPacket_f_reg[7][30]  ( .CLK(n5929), .D(N10608), .Q(
        decodedPacket7_o[30]) );
  LATCHX1 \decodedPacket_f_reg[7][29]  ( .CLK(n5929), .D(N10607), .Q(
        decodedPacket7_o[29]) );
  LATCHX1 \decodedPacket_f_reg[7][28]  ( .CLK(n5929), .D(N10606), .Q(
        decodedPacket7_o[28]) );
  LATCHX1 \decodedPacket_f_reg[7][27]  ( .CLK(n5929), .D(N10605), .Q(
        decodedPacket7_o[27]) );
  LATCHX1 \decodedPacket_f_reg[7][26]  ( .CLK(n5929), .D(N10604), .Q(
        decodedPacket7_o[26]) );
  LATCHX1 \decodedPacket_f_reg[7][25]  ( .CLK(n5929), .D(N10603), .Q(
        decodedPacket7_o[25]) );
  LATCHX1 \decodedPacket_f_reg[7][24]  ( .CLK(n5929), .D(N10602), .Q(
        decodedPacket7_o[24]) );
  LATCHX1 \decodedPacket_f_reg[7][23]  ( .CLK(n5928), .D(N10601), .Q(
        decodedPacket7_o[23]) );
  LATCHX1 \decodedPacket_f_reg[7][22]  ( .CLK(n5928), .D(N10600), .Q(
        decodedPacket7_o[22]) );
  LATCHX1 \decodedPacket_f_reg[7][21]  ( .CLK(n5928), .D(N10599), .Q(
        decodedPacket7_o[21]) );
  LATCHX1 \decodedPacket_f_reg[7][20]  ( .CLK(n5928), .D(N10598), .Q(
        decodedPacket7_o[20]) );
  LATCHX1 \decodedPacket_f_reg[7][19]  ( .CLK(n5928), .D(N10597), .Q(
        decodedPacket7_o[19]) );
  LATCHX1 \decodedPacket_f_reg[7][18]  ( .CLK(n5928), .D(N10596), .Q(
        decodedPacket7_o[18]) );
  LATCHX1 \decodedPacket_f_reg[7][17]  ( .CLK(n5928), .D(N10595), .Q(
        decodedPacket7_o[17]) );
  LATCHX1 \decodedPacket_f_reg[7][16]  ( .CLK(n5928), .D(N10594), .Q(
        decodedPacket7_o[16]) );
  LATCHX1 \decodedPacket_f_reg[7][15]  ( .CLK(n5928), .D(N10593), .Q(
        decodedPacket7_o[15]) );
  LATCHX1 \decodedPacket_f_reg[7][14]  ( .CLK(n5928), .D(N10592), .Q(
        decodedPacket7_o[14]) );
  LATCHX1 \decodedPacket_f_reg[7][13]  ( .CLK(n5928), .D(N10591), .Q(
        decodedPacket7_o[13]) );
  LATCHX1 \decodedPacket_f_reg[7][12]  ( .CLK(n5928), .D(N10590), .Q(
        decodedPacket7_o[12]) );
  LATCHX1 \decodedPacket_f_reg[7][11]  ( .CLK(n5927), .D(N10589), .Q(
        decodedPacket7_o[11]) );
  LATCHX1 \decodedPacket_f_reg[7][10]  ( .CLK(n5927), .D(N10588), .Q(
        decodedPacket7_o[10]) );
  LATCHX1 \decodedPacket_f_reg[7][9]  ( .CLK(n5927), .D(N10587), .Q(
        decodedPacket7_o[9]) );
  LATCHX1 \decodedPacket_f_reg[7][8]  ( .CLK(n5927), .D(N10586), .Q(
        decodedPacket7_o[8]) );
  LATCHX1 \decodedPacket_f_reg[7][7]  ( .CLK(n5927), .D(N10585), .Q(
        decodedPacket7_o[7]) );
  LATCHX1 \decodedPacket_f_reg[7][6]  ( .CLK(n5927), .D(N10584), .Q(
        decodedPacket7_o[6]) );
  LATCHX1 \decodedPacket_f_reg[7][5]  ( .CLK(n5927), .D(N10583), .Q(
        decodedPacket7_o[5]) );
  LATCHX1 \decodedPacket_f_reg[7][4]  ( .CLK(n5927), .D(N10582), .Q(
        decodedPacket7_o[4]) );
  LATCHX1 \decodedPacket_f_reg[7][3]  ( .CLK(n5927), .D(N10581), .Q(
        decodedPacket7_o[3]) );
  LATCHX1 \decodedPacket_f_reg[7][2]  ( .CLK(n5927), .D(N10580), .Q(
        decodedPacket7_o[2]) );
  LATCHX1 \decodedPacket_f_reg[7][1]  ( .CLK(n5927), .D(N10579), .Q(
        decodedPacket7_o[1]) );
  LATCHX1 \decodedPacket_f_reg[7][0]  ( .CLK(n5927), .D(N10578), .Q(
        decodedPacket7_o[0]) );
  LATCHX1 \decodedPacket_f_reg[6][121]  ( .CLK(n5921), .D(N10572), .Q(
        decodedPacket6_o[121]) );
  LATCHX1 \decodedPacket_f_reg[6][120]  ( .CLK(n5922), .D(N10571), .Q(
        decodedPacket6_o[120]) );
  LATCHX1 \decodedPacket_f_reg[6][119]  ( .CLK(n5926), .D(N10570), .Q(
        decodedPacket6_o[119]) );
  LATCHX1 \decodedPacket_f_reg[6][118]  ( .CLK(n5926), .D(N10569), .Q(
        decodedPacket6_o[118]) );
  LATCHX1 \decodedPacket_f_reg[6][117]  ( .CLK(n5926), .D(N10568), .Q(
        decodedPacket6_o[117]) );
  LATCHX1 \decodedPacket_f_reg[6][116]  ( .CLK(n5926), .D(N10567), .Q(
        decodedPacket6_o[116]) );
  LATCHX1 \decodedPacket_f_reg[6][115]  ( .CLK(n5926), .D(N10566), .Q(
        decodedPacket6_o[115]) );
  LATCHX1 \decodedPacket_f_reg[6][114]  ( .CLK(n5926), .D(N10565), .Q(
        decodedPacket6_o[114]) );
  LATCHX1 \decodedPacket_f_reg[6][113]  ( .CLK(n5926), .D(N10564), .Q(
        decodedPacket6_o[113]) );
  LATCHX1 \decodedPacket_f_reg[6][112]  ( .CLK(n5926), .D(N10563), .Q(
        decodedPacket6_o[112]) );
  LATCHX1 \decodedPacket_f_reg[6][111]  ( .CLK(n5926), .D(N10562), .Q(
        decodedPacket6_o[111]) );
  LATCHX1 \decodedPacket_f_reg[6][110]  ( .CLK(n5926), .D(N10561), .Q(
        decodedPacket6_o[110]) );
  LATCHX1 \decodedPacket_f_reg[6][109]  ( .CLK(n5926), .D(N10560), .Q(
        decodedPacket6_o[109]) );
  LATCHX1 \decodedPacket_f_reg[6][108]  ( .CLK(n5926), .D(N10559), .Q(
        decodedPacket6_o[108]) );
  LATCHX1 \decodedPacket_f_reg[6][107]  ( .CLK(n5925), .D(N10558), .Q(
        decodedPacket6_o[107]) );
  LATCHX1 \decodedPacket_f_reg[6][106]  ( .CLK(n5925), .D(N10557), .Q(
        decodedPacket6_o[106]) );
  LATCHX1 \decodedPacket_f_reg[6][105]  ( .CLK(n5925), .D(N10556), .Q(
        decodedPacket6_o[105]) );
  LATCHX1 \decodedPacket_f_reg[6][104]  ( .CLK(n5925), .D(N10555), .Q(
        decodedPacket6_o[104]) );
  LATCHX1 \decodedPacket_f_reg[6][103]  ( .CLK(n5925), .D(N10554), .Q(
        decodedPacket6_o[103]) );
  LATCHX1 \decodedPacket_f_reg[6][102]  ( .CLK(n5925), .D(N10553), .Q(
        decodedPacket6_o[102]) );
  LATCHX1 \decodedPacket_f_reg[6][101]  ( .CLK(n5925), .D(N10552), .Q(
        decodedPacket6_o[101]) );
  LATCHX1 \decodedPacket_f_reg[6][100]  ( .CLK(n5925), .D(N10551), .Q(
        decodedPacket6_o[100]) );
  LATCHX1 \decodedPacket_f_reg[6][99]  ( .CLK(n5925), .D(N10550), .Q(
        decodedPacket6_o[99]) );
  LATCHX1 \decodedPacket_f_reg[6][98]  ( .CLK(n5925), .D(N10548), .Q(
        decodedPacket6_o[98]) );
  LATCHX1 \decodedPacket_f_reg[6][97]  ( .CLK(n5925), .D(N10546), .Q(
        decodedPacket6_o[97]) );
  LATCHX1 \decodedPacket_f_reg[6][96]  ( .CLK(n5925), .D(N10545), .Q(
        decodedPacket6_o[96]) );
  LATCHX1 \decodedPacket_f_reg[6][95]  ( .CLK(n5924), .D(N10544), .Q(
        decodedPacket6_o[95]) );
  LATCHX1 \decodedPacket_f_reg[6][94]  ( .CLK(n5924), .D(N10543), .Q(
        decodedPacket6_o[94]) );
  LATCHX1 \decodedPacket_f_reg[6][93]  ( .CLK(n5924), .D(N10542), .Q(
        decodedPacket6_o[93]) );
  LATCHX1 \decodedPacket_f_reg[6][92]  ( .CLK(n5924), .D(N10541), .Q(
        decodedPacket6_o[92]) );
  LATCHX1 \decodedPacket_f_reg[6][91]  ( .CLK(n5924), .D(N10540), .Q(
        decodedPacket6_o[91]) );
  LATCHX1 \decodedPacket_f_reg[6][90]  ( .CLK(n5924), .D(N10539), .Q(
        decodedPacket6_o[90]) );
  LATCHX1 \decodedPacket_f_reg[6][89]  ( .CLK(n5924), .D(N10538), .Q(
        decodedPacket6_o[89]) );
  LATCHX1 \decodedPacket_f_reg[6][88]  ( .CLK(n5924), .D(N10537), .Q(
        decodedPacket6_o[88]) );
  LATCHX1 \decodedPacket_f_reg[6][87]  ( .CLK(n5924), .D(N10536), .Q(
        decodedPacket6_o[87]) );
  LATCHX1 \decodedPacket_f_reg[6][86]  ( .CLK(n5924), .D(N10535), .Q(
        decodedPacket6_o[86]) );
  LATCHX1 \decodedPacket_f_reg[6][85]  ( .CLK(n5924), .D(N10534), .Q(
        decodedPacket6_o[85]) );
  LATCHX1 \decodedPacket_f_reg[6][84]  ( .CLK(n5924), .D(N10533), .Q(
        decodedPacket6_o[84]) );
  LATCHX1 \decodedPacket_f_reg[6][83]  ( .CLK(n5923), .D(N10532), .Q(
        decodedPacket6_o[83]) );
  LATCHX1 \decodedPacket_f_reg[6][82]  ( .CLK(n5923), .D(N10531), .Q(
        decodedPacket6_o[82]) );
  LATCHX1 \decodedPacket_f_reg[6][81]  ( .CLK(n5923), .D(N10530), .Q(
        decodedPacket6_o[81]) );
  LATCHX1 \decodedPacket_f_reg[6][80]  ( .CLK(n5923), .D(N10529), .Q(
        decodedPacket6_o[80]) );
  LATCHX1 \decodedPacket_f_reg[6][79]  ( .CLK(n5923), .D(N10528), .Q(
        decodedPacket6_o[79]) );
  LATCHX1 \decodedPacket_f_reg[6][78]  ( .CLK(n5923), .D(N10527), .Q(
        decodedPacket6_o[78]) );
  LATCHX1 \decodedPacket_f_reg[6][77]  ( .CLK(n5923), .D(N10526), .Q(
        decodedPacket6_o[77]) );
  LATCHX1 \decodedPacket_f_reg[6][76]  ( .CLK(n5923), .D(N10525), .Q(
        decodedPacket6_o[76]) );
  LATCHX1 \decodedPacket_f_reg[6][75]  ( .CLK(n5923), .D(N10524), .Q(
        decodedPacket6_o[75]) );
  LATCHX1 \decodedPacket_f_reg[6][74]  ( .CLK(n5923), .D(N10523), .Q(
        decodedPacket6_o[74]) );
  LATCHX1 \decodedPacket_f_reg[6][73]  ( .CLK(n5923), .D(N10522), .Q(
        decodedPacket6_o[73]) );
  LATCHX1 \decodedPacket_f_reg[6][72]  ( .CLK(n5923), .D(N10521), .Q(
        decodedPacket6_o[72]) );
  LATCHX1 \decodedPacket_f_reg[6][71]  ( .CLK(n5922), .D(N10520), .Q(
        decodedPacket6_o[71]) );
  LATCHX1 \decodedPacket_f_reg[6][70]  ( .CLK(n5922), .D(N10519), .Q(
        decodedPacket6_o[70]) );
  LATCHX1 \decodedPacket_f_reg[6][69]  ( .CLK(n5922), .D(N10518), .Q(
        decodedPacket6_o[69]) );
  LATCHX1 \decodedPacket_f_reg[6][68]  ( .CLK(n5922), .D(N10517), .Q(
        decodedPacket6_o[68]) );
  LATCHX1 \decodedPacket_f_reg[6][67]  ( .CLK(n5922), .D(N10516), .Q(
        decodedPacket6_o[67]) );
  LATCHX1 \decodedPacket_f_reg[6][66]  ( .CLK(n5922), .D(N10515), .Q(
        decodedPacket6_o[66]) );
  LATCHX1 \decodedPacket_f_reg[6][65]  ( .CLK(n5922), .D(N10514), .Q(
        decodedPacket6_o[65]) );
  LATCHX1 \decodedPacket_f_reg[6][64]  ( .CLK(n5922), .D(N10513), .Q(
        decodedPacket6_o[64]) );
  LATCHX1 \decodedPacket_f_reg[6][63]  ( .CLK(n5922), .D(N10512), .Q(
        decodedPacket6_o[63]) );
  LATCHX1 \decodedPacket_f_reg[6][62]  ( .CLK(n5922), .D(N10511), .Q(
        decodedPacket6_o[62]) );
  LATCHX1 \decodedPacket_f_reg[6][61]  ( .CLK(n5922), .D(N10510), .Q(
        decodedPacket6_o[61]) );
  LATCHX1 \decodedPacket_f_reg[6][60]  ( .CLK(n5922), .D(N10509), .Q(
        decodedPacket6_o[60]) );
  LATCHX1 \decodedPacket_f_reg[6][59]  ( .CLK(n5921), .D(N10508), .Q(
        decodedPacket6_o[59]) );
  LATCHX1 \decodedPacket_f_reg[6][58]  ( .CLK(n5921), .D(N10507), .Q(
        decodedPacket6_o[58]) );
  LATCHX1 \decodedPacket_f_reg[6][57]  ( .CLK(n5921), .D(N10506), .Q(
        decodedPacket6_o[57]) );
  LATCHX1 \decodedPacket_f_reg[6][56]  ( .CLK(n5921), .D(N10505), .Q(
        decodedPacket6_o[56]) );
  LATCHX1 \decodedPacket_f_reg[6][55]  ( .CLK(n5921), .D(N10504), .Q(
        decodedPacket6_o[55]) );
  LATCHX1 \decodedPacket_f_reg[6][54]  ( .CLK(n5921), .D(N10503), .Q(
        decodedPacket6_o[54]) );
  LATCHX1 \decodedPacket_f_reg[6][53]  ( .CLK(n5921), .D(N10502), .Q(
        decodedPacket6_o[53]) );
  LATCHX1 \decodedPacket_f_reg[6][52]  ( .CLK(n5921), .D(N10501), .Q(
        decodedPacket6_o[52]) );
  LATCHX1 \decodedPacket_f_reg[6][51]  ( .CLK(n5921), .D(N10500), .Q(
        decodedPacket6_o[51]) );
  LATCHX1 \decodedPacket_f_reg[6][50]  ( .CLK(n5921), .D(N10499), .Q(
        decodedPacket6_o[50]) );
  LATCHX1 \decodedPacket_f_reg[6][49]  ( .CLK(n5921), .D(N10498), .Q(
        decodedPacket6_o[49]) );
  LATCHX1 \decodedPacket_f_reg[6][48]  ( .CLK(n5921), .D(N10496), .Q(
        decodedPacket6_o[48]) );
  LATCHX1 \decodedPacket_f_reg[6][47]  ( .CLK(n5920), .D(N10495), .Q(
        decodedPacket6_o[47]) );
  LATCHX1 \decodedPacket_f_reg[6][46]  ( .CLK(n5920), .D(N10494), .Q(
        decodedPacket6_o[46]) );
  LATCHX1 \decodedPacket_f_reg[6][45]  ( .CLK(n5920), .D(N10493), .Q(
        decodedPacket6_o[45]) );
  LATCHX1 \decodedPacket_f_reg[6][44]  ( .CLK(n5920), .D(N10492), .Q(
        decodedPacket6_o[44]) );
  LATCHX1 \decodedPacket_f_reg[6][43]  ( .CLK(n5920), .D(N10491), .Q(
        decodedPacket6_o[43]) );
  LATCHX1 \decodedPacket_f_reg[6][42]  ( .CLK(n5920), .D(N10490), .Q(
        decodedPacket6_o[42]) );
  LATCHX1 \decodedPacket_f_reg[6][41]  ( .CLK(n5920), .D(N10489), .Q(
        decodedPacket6_o[41]) );
  LATCHX1 \decodedPacket_f_reg[6][40]  ( .CLK(n5920), .D(N10488), .Q(
        decodedPacket6_o[40]) );
  LATCHX1 \decodedPacket_f_reg[6][39]  ( .CLK(n5920), .D(N10487), .Q(
        decodedPacket6_o[39]) );
  LATCHX1 \decodedPacket_f_reg[6][38]  ( .CLK(n5920), .D(N10486), .Q(
        decodedPacket6_o[38]) );
  LATCHX1 \decodedPacket_f_reg[6][37]  ( .CLK(n5920), .D(N10485), .Q(
        decodedPacket6_o[37]) );
  LATCHX1 \decodedPacket_f_reg[6][36]  ( .CLK(n5920), .D(N10484), .Q(
        decodedPacket6_o[36]) );
  LATCHX1 \decodedPacket_f_reg[6][35]  ( .CLK(n5919), .D(N10483), .Q(
        decodedPacket6_o[35]) );
  LATCHX1 \decodedPacket_f_reg[6][34]  ( .CLK(n5919), .D(N10482), .Q(
        decodedPacket6_o[34]) );
  LATCHX1 \decodedPacket_f_reg[6][33]  ( .CLK(n5919), .D(N10481), .Q(
        decodedPacket6_o[33]) );
  LATCHX1 \decodedPacket_f_reg[6][32]  ( .CLK(n5919), .D(N10480), .Q(
        decodedPacket6_o[32]) );
  LATCHX1 \decodedPacket_f_reg[6][31]  ( .CLK(n5919), .D(N10479), .Q(
        decodedPacket6_o[31]) );
  LATCHX1 \decodedPacket_f_reg[6][30]  ( .CLK(n5919), .D(N10478), .Q(
        decodedPacket6_o[30]) );
  LATCHX1 \decodedPacket_f_reg[6][29]  ( .CLK(n5919), .D(N10477), .Q(
        decodedPacket6_o[29]) );
  LATCHX1 \decodedPacket_f_reg[6][28]  ( .CLK(n5919), .D(N10476), .Q(
        decodedPacket6_o[28]) );
  LATCHX1 \decodedPacket_f_reg[6][27]  ( .CLK(n5919), .D(N10475), .Q(
        decodedPacket6_o[27]) );
  LATCHX1 \decodedPacket_f_reg[6][26]  ( .CLK(n5919), .D(N10474), .Q(
        decodedPacket6_o[26]) );
  LATCHX1 \decodedPacket_f_reg[6][25]  ( .CLK(n5919), .D(N10473), .Q(
        decodedPacket6_o[25]) );
  LATCHX1 \decodedPacket_f_reg[6][24]  ( .CLK(n5919), .D(N10472), .Q(
        decodedPacket6_o[24]) );
  LATCHX1 \decodedPacket_f_reg[6][23]  ( .CLK(n5918), .D(N10471), .Q(
        decodedPacket6_o[23]) );
  LATCHX1 \decodedPacket_f_reg[6][22]  ( .CLK(n5918), .D(N10470), .Q(
        decodedPacket6_o[22]) );
  LATCHX1 \decodedPacket_f_reg[6][21]  ( .CLK(n5918), .D(N10469), .Q(
        decodedPacket6_o[21]) );
  LATCHX1 \decodedPacket_f_reg[6][20]  ( .CLK(n5918), .D(N10468), .Q(
        decodedPacket6_o[20]) );
  LATCHX1 \decodedPacket_f_reg[6][19]  ( .CLK(n5918), .D(N10467), .Q(
        decodedPacket6_o[19]) );
  LATCHX1 \decodedPacket_f_reg[6][18]  ( .CLK(n5918), .D(N10466), .Q(
        decodedPacket6_o[18]) );
  LATCHX1 \decodedPacket_f_reg[6][17]  ( .CLK(n5918), .D(N10465), .Q(
        decodedPacket6_o[17]) );
  LATCHX1 \decodedPacket_f_reg[6][16]  ( .CLK(n5918), .D(N10464), .Q(
        decodedPacket6_o[16]) );
  LATCHX1 \decodedPacket_f_reg[6][15]  ( .CLK(n5918), .D(N10463), .Q(
        decodedPacket6_o[15]) );
  LATCHX1 \decodedPacket_f_reg[6][14]  ( .CLK(n5918), .D(N10462), .Q(
        decodedPacket6_o[14]) );
  LATCHX1 \decodedPacket_f_reg[6][13]  ( .CLK(n5918), .D(N10461), .Q(
        decodedPacket6_o[13]) );
  LATCHX1 \decodedPacket_f_reg[6][12]  ( .CLK(n5918), .D(N10460), .Q(
        decodedPacket6_o[12]) );
  LATCHX1 \decodedPacket_f_reg[6][11]  ( .CLK(n5917), .D(N10459), .Q(
        decodedPacket6_o[11]) );
  LATCHX1 \decodedPacket_f_reg[6][10]  ( .CLK(n5917), .D(N10458), .Q(
        decodedPacket6_o[10]) );
  LATCHX1 \decodedPacket_f_reg[6][9]  ( .CLK(n5917), .D(N10457), .Q(
        decodedPacket6_o[9]) );
  LATCHX1 \decodedPacket_f_reg[6][8]  ( .CLK(n5917), .D(N10456), .Q(
        decodedPacket6_o[8]) );
  LATCHX1 \decodedPacket_f_reg[6][7]  ( .CLK(n5917), .D(N10455), .Q(
        decodedPacket6_o[7]) );
  LATCHX1 \decodedPacket_f_reg[6][6]  ( .CLK(n5917), .D(N10454), .Q(
        decodedPacket6_o[6]) );
  LATCHX1 \decodedPacket_f_reg[6][5]  ( .CLK(n5917), .D(N10453), .Q(
        decodedPacket6_o[5]) );
  LATCHX1 \decodedPacket_f_reg[6][4]  ( .CLK(n5917), .D(N10452), .Q(
        decodedPacket6_o[4]) );
  LATCHX1 \decodedPacket_f_reg[6][3]  ( .CLK(n5917), .D(N10451), .Q(
        decodedPacket6_o[3]) );
  LATCHX1 \decodedPacket_f_reg[6][2]  ( .CLK(n5917), .D(N10450), .Q(
        decodedPacket6_o[2]) );
  LATCHX1 \decodedPacket_f_reg[6][1]  ( .CLK(n5917), .D(N10449), .Q(
        decodedPacket6_o[1]) );
  LATCHX1 \decodedPacket_f_reg[6][0]  ( .CLK(n5917), .D(N10448), .Q(
        decodedPacket6_o[0]) );
  LATCHX1 \decodedPacket_f_reg[5][121]  ( .CLK(n5911), .D(N10442), .Q(
        decodedPacket5_o[121]) );
  LATCHX1 \decodedPacket_f_reg[5][120]  ( .CLK(n5912), .D(N10441), .Q(
        decodedPacket5_o[120]) );
  LATCHX1 \decodedPacket_f_reg[5][119]  ( .CLK(n5916), .D(N10440), .Q(
        decodedPacket5_o[119]) );
  LATCHX1 \decodedPacket_f_reg[5][118]  ( .CLK(n5916), .D(N10439), .Q(
        decodedPacket5_o[118]) );
  LATCHX1 \decodedPacket_f_reg[5][117]  ( .CLK(n5916), .D(N10438), .Q(
        decodedPacket5_o[117]) );
  LATCHX1 \decodedPacket_f_reg[5][116]  ( .CLK(n5916), .D(N10437), .Q(
        decodedPacket5_o[116]) );
  LATCHX1 \decodedPacket_f_reg[5][115]  ( .CLK(n5916), .D(N10436), .Q(
        decodedPacket5_o[115]) );
  LATCHX1 \decodedPacket_f_reg[5][114]  ( .CLK(n5916), .D(N10435), .Q(
        decodedPacket5_o[114]) );
  LATCHX1 \decodedPacket_f_reg[5][113]  ( .CLK(n5916), .D(N10434), .Q(
        decodedPacket5_o[113]) );
  LATCHX1 \decodedPacket_f_reg[5][112]  ( .CLK(n5916), .D(N10433), .Q(
        decodedPacket5_o[112]) );
  LATCHX1 \decodedPacket_f_reg[5][111]  ( .CLK(n5916), .D(N10432), .Q(
        decodedPacket5_o[111]) );
  LATCHX1 \decodedPacket_f_reg[5][110]  ( .CLK(n5916), .D(N10431), .Q(
        decodedPacket5_o[110]) );
  LATCHX1 \decodedPacket_f_reg[5][109]  ( .CLK(n5916), .D(N10430), .Q(
        decodedPacket5_o[109]) );
  LATCHX1 \decodedPacket_f_reg[5][108]  ( .CLK(n5916), .D(N10429), .Q(
        decodedPacket5_o[108]) );
  LATCHX1 \decodedPacket_f_reg[5][107]  ( .CLK(n5915), .D(N10428), .Q(
        decodedPacket5_o[107]) );
  LATCHX1 \decodedPacket_f_reg[5][106]  ( .CLK(n5915), .D(N10427), .Q(
        decodedPacket5_o[106]) );
  LATCHX1 \decodedPacket_f_reg[5][105]  ( .CLK(n5915), .D(N10426), .Q(
        decodedPacket5_o[105]) );
  LATCHX1 \decodedPacket_f_reg[5][104]  ( .CLK(n5915), .D(N10425), .Q(
        decodedPacket5_o[104]) );
  LATCHX1 \decodedPacket_f_reg[5][103]  ( .CLK(n5915), .D(N10424), .Q(
        decodedPacket5_o[103]) );
  LATCHX1 \decodedPacket_f_reg[5][102]  ( .CLK(n5915), .D(N10423), .Q(
        decodedPacket5_o[102]) );
  LATCHX1 \decodedPacket_f_reg[5][101]  ( .CLK(n5915), .D(N10422), .Q(
        decodedPacket5_o[101]) );
  LATCHX1 \decodedPacket_f_reg[5][100]  ( .CLK(n5915), .D(N10421), .Q(
        decodedPacket5_o[100]) );
  LATCHX1 \decodedPacket_f_reg[5][99]  ( .CLK(n5915), .D(N10420), .Q(
        decodedPacket5_o[99]) );
  LATCHX1 \decodedPacket_f_reg[5][98]  ( .CLK(n5915), .D(N10418), .Q(
        decodedPacket5_o[98]) );
  LATCHX1 \decodedPacket_f_reg[5][97]  ( .CLK(n5915), .D(N10416), .Q(
        decodedPacket5_o[97]) );
  LATCHX1 \decodedPacket_f_reg[5][96]  ( .CLK(n5915), .D(N10415), .Q(
        decodedPacket5_o[96]) );
  LATCHX1 \decodedPacket_f_reg[5][95]  ( .CLK(n5914), .D(N10414), .Q(
        decodedPacket5_o[95]) );
  LATCHX1 \decodedPacket_f_reg[5][94]  ( .CLK(n5914), .D(N10413), .Q(
        decodedPacket5_o[94]) );
  LATCHX1 \decodedPacket_f_reg[5][93]  ( .CLK(n5914), .D(N10412), .Q(
        decodedPacket5_o[93]) );
  LATCHX1 \decodedPacket_f_reg[5][92]  ( .CLK(n5914), .D(N10411), .Q(
        decodedPacket5_o[92]) );
  LATCHX1 \decodedPacket_f_reg[5][91]  ( .CLK(n5914), .D(N10410), .Q(
        decodedPacket5_o[91]) );
  LATCHX1 \decodedPacket_f_reg[5][90]  ( .CLK(n5914), .D(N10409), .Q(
        decodedPacket5_o[90]) );
  LATCHX1 \decodedPacket_f_reg[5][89]  ( .CLK(n5914), .D(N10408), .Q(
        decodedPacket5_o[89]) );
  LATCHX1 \decodedPacket_f_reg[5][88]  ( .CLK(n5914), .D(N10407), .Q(
        decodedPacket5_o[88]) );
  LATCHX1 \decodedPacket_f_reg[5][87]  ( .CLK(n5914), .D(N10406), .Q(
        decodedPacket5_o[87]) );
  LATCHX1 \decodedPacket_f_reg[5][86]  ( .CLK(n5914), .D(N10405), .Q(
        decodedPacket5_o[86]) );
  LATCHX1 \decodedPacket_f_reg[5][85]  ( .CLK(n5914), .D(N10404), .Q(
        decodedPacket5_o[85]) );
  LATCHX1 \decodedPacket_f_reg[5][84]  ( .CLK(n5914), .D(N10403), .Q(
        decodedPacket5_o[84]) );
  LATCHX1 \decodedPacket_f_reg[5][83]  ( .CLK(n5913), .D(N10402), .Q(
        decodedPacket5_o[83]) );
  LATCHX1 \decodedPacket_f_reg[5][82]  ( .CLK(n5913), .D(N10401), .Q(
        decodedPacket5_o[82]) );
  LATCHX1 \decodedPacket_f_reg[5][81]  ( .CLK(n5913), .D(N10400), .Q(
        decodedPacket5_o[81]) );
  LATCHX1 \decodedPacket_f_reg[5][80]  ( .CLK(n5913), .D(N10399), .Q(
        decodedPacket5_o[80]) );
  LATCHX1 \decodedPacket_f_reg[5][79]  ( .CLK(n5913), .D(N10398), .Q(
        decodedPacket5_o[79]) );
  LATCHX1 \decodedPacket_f_reg[5][78]  ( .CLK(n5913), .D(N10397), .Q(
        decodedPacket5_o[78]) );
  LATCHX1 \decodedPacket_f_reg[5][77]  ( .CLK(n5913), .D(N10396), .Q(
        decodedPacket5_o[77]) );
  LATCHX1 \decodedPacket_f_reg[5][76]  ( .CLK(n5913), .D(N10395), .Q(
        decodedPacket5_o[76]) );
  LATCHX1 \decodedPacket_f_reg[5][75]  ( .CLK(n5913), .D(N10394), .Q(
        decodedPacket5_o[75]) );
  LATCHX1 \decodedPacket_f_reg[5][74]  ( .CLK(n5913), .D(N10393), .Q(
        decodedPacket5_o[74]) );
  LATCHX1 \decodedPacket_f_reg[5][73]  ( .CLK(n5913), .D(N10392), .Q(
        decodedPacket5_o[73]) );
  LATCHX1 \decodedPacket_f_reg[5][72]  ( .CLK(n5913), .D(N10391), .Q(
        decodedPacket5_o[72]) );
  LATCHX1 \decodedPacket_f_reg[5][71]  ( .CLK(n5912), .D(N10390), .Q(
        decodedPacket5_o[71]) );
  LATCHX1 \decodedPacket_f_reg[5][70]  ( .CLK(n5912), .D(N10389), .Q(
        decodedPacket5_o[70]) );
  LATCHX1 \decodedPacket_f_reg[5][69]  ( .CLK(n5912), .D(N10388), .Q(
        decodedPacket5_o[69]) );
  LATCHX1 \decodedPacket_f_reg[5][68]  ( .CLK(n5912), .D(N10387), .Q(
        decodedPacket5_o[68]) );
  LATCHX1 \decodedPacket_f_reg[5][67]  ( .CLK(n5912), .D(N10386), .Q(
        decodedPacket5_o[67]) );
  LATCHX1 \decodedPacket_f_reg[5][66]  ( .CLK(n5912), .D(N10385), .Q(
        decodedPacket5_o[66]) );
  LATCHX1 \decodedPacket_f_reg[5][65]  ( .CLK(n5912), .D(N10384), .Q(
        decodedPacket5_o[65]) );
  LATCHX1 \decodedPacket_f_reg[5][64]  ( .CLK(n5912), .D(N10383), .Q(
        decodedPacket5_o[64]) );
  LATCHX1 \decodedPacket_f_reg[5][63]  ( .CLK(n5912), .D(N10382), .Q(
        decodedPacket5_o[63]) );
  LATCHX1 \decodedPacket_f_reg[5][62]  ( .CLK(n5912), .D(N10381), .Q(
        decodedPacket5_o[62]) );
  LATCHX1 \decodedPacket_f_reg[5][61]  ( .CLK(n5912), .D(N10380), .Q(
        decodedPacket5_o[61]) );
  LATCHX1 \decodedPacket_f_reg[5][60]  ( .CLK(n5912), .D(N10379), .Q(
        decodedPacket5_o[60]) );
  LATCHX1 \decodedPacket_f_reg[5][59]  ( .CLK(n5911), .D(N10378), .Q(
        decodedPacket5_o[59]) );
  LATCHX1 \decodedPacket_f_reg[5][58]  ( .CLK(n5911), .D(N10377), .Q(
        decodedPacket5_o[58]) );
  LATCHX1 \decodedPacket_f_reg[5][57]  ( .CLK(n5911), .D(N10376), .Q(
        decodedPacket5_o[57]) );
  LATCHX1 \decodedPacket_f_reg[5][56]  ( .CLK(n5911), .D(N10375), .Q(
        decodedPacket5_o[56]) );
  LATCHX1 \decodedPacket_f_reg[5][55]  ( .CLK(n5911), .D(N10374), .Q(
        decodedPacket5_o[55]) );
  LATCHX1 \decodedPacket_f_reg[5][54]  ( .CLK(n5911), .D(N10373), .Q(
        decodedPacket5_o[54]) );
  LATCHX1 \decodedPacket_f_reg[5][53]  ( .CLK(n5911), .D(N10372), .Q(
        decodedPacket5_o[53]) );
  LATCHX1 \decodedPacket_f_reg[5][52]  ( .CLK(n5911), .D(N10371), .Q(
        decodedPacket5_o[52]) );
  LATCHX1 \decodedPacket_f_reg[5][51]  ( .CLK(n5911), .D(N10370), .Q(
        decodedPacket5_o[51]) );
  LATCHX1 \decodedPacket_f_reg[5][50]  ( .CLK(n5911), .D(N10369), .Q(
        decodedPacket5_o[50]) );
  LATCHX1 \decodedPacket_f_reg[5][49]  ( .CLK(n5911), .D(N10368), .Q(
        decodedPacket5_o[49]) );
  LATCHX1 \decodedPacket_f_reg[5][48]  ( .CLK(n5911), .D(N10366), .Q(
        decodedPacket5_o[48]) );
  LATCHX1 \decodedPacket_f_reg[5][47]  ( .CLK(n5910), .D(N10365), .Q(
        decodedPacket5_o[47]) );
  LATCHX1 \decodedPacket_f_reg[5][46]  ( .CLK(n5910), .D(N10364), .Q(
        decodedPacket5_o[46]) );
  LATCHX1 \decodedPacket_f_reg[5][45]  ( .CLK(n5910), .D(N10363), .Q(
        decodedPacket5_o[45]) );
  LATCHX1 \decodedPacket_f_reg[5][44]  ( .CLK(n5910), .D(N10362), .Q(
        decodedPacket5_o[44]) );
  LATCHX1 \decodedPacket_f_reg[5][43]  ( .CLK(n5910), .D(N10361), .Q(
        decodedPacket5_o[43]) );
  LATCHX1 \decodedPacket_f_reg[5][42]  ( .CLK(n5910), .D(N10360), .Q(
        decodedPacket5_o[42]) );
  LATCHX1 \decodedPacket_f_reg[5][41]  ( .CLK(n5910), .D(N10359), .Q(
        decodedPacket5_o[41]) );
  LATCHX1 \decodedPacket_f_reg[5][40]  ( .CLK(n5910), .D(N10358), .Q(
        decodedPacket5_o[40]) );
  LATCHX1 \decodedPacket_f_reg[5][39]  ( .CLK(n5910), .D(N10357), .Q(
        decodedPacket5_o[39]) );
  LATCHX1 \decodedPacket_f_reg[5][38]  ( .CLK(n5910), .D(N10356), .Q(
        decodedPacket5_o[38]) );
  LATCHX1 \decodedPacket_f_reg[5][37]  ( .CLK(n5910), .D(N10355), .Q(
        decodedPacket5_o[37]) );
  LATCHX1 \decodedPacket_f_reg[5][36]  ( .CLK(n5910), .D(N10354), .Q(
        decodedPacket5_o[36]) );
  LATCHX1 \decodedPacket_f_reg[5][35]  ( .CLK(n5909), .D(N10353), .Q(
        decodedPacket5_o[35]) );
  LATCHX1 \decodedPacket_f_reg[5][34]  ( .CLK(n5909), .D(N10352), .Q(
        decodedPacket5_o[34]) );
  LATCHX1 \decodedPacket_f_reg[5][33]  ( .CLK(n5909), .D(N10351), .Q(
        decodedPacket5_o[33]) );
  LATCHX1 \decodedPacket_f_reg[5][32]  ( .CLK(n5909), .D(N10350), .Q(
        decodedPacket5_o[32]) );
  LATCHX1 \decodedPacket_f_reg[5][31]  ( .CLK(n5909), .D(N10349), .Q(
        decodedPacket5_o[31]) );
  LATCHX1 \decodedPacket_f_reg[5][30]  ( .CLK(n5909), .D(N10348), .Q(
        decodedPacket5_o[30]) );
  LATCHX1 \decodedPacket_f_reg[5][29]  ( .CLK(n5909), .D(N10347), .Q(
        decodedPacket5_o[29]) );
  LATCHX1 \decodedPacket_f_reg[5][28]  ( .CLK(n5909), .D(N10346), .Q(
        decodedPacket5_o[28]) );
  LATCHX1 \decodedPacket_f_reg[5][27]  ( .CLK(n5909), .D(N10345), .Q(
        decodedPacket5_o[27]) );
  LATCHX1 \decodedPacket_f_reg[5][26]  ( .CLK(n5909), .D(N10344), .Q(
        decodedPacket5_o[26]) );
  LATCHX1 \decodedPacket_f_reg[5][25]  ( .CLK(n5909), .D(N10343), .Q(
        decodedPacket5_o[25]) );
  LATCHX1 \decodedPacket_f_reg[5][24]  ( .CLK(n5909), .D(N10342), .Q(
        decodedPacket5_o[24]) );
  LATCHX1 \decodedPacket_f_reg[5][23]  ( .CLK(n5908), .D(N10341), .Q(
        decodedPacket5_o[23]) );
  LATCHX1 \decodedPacket_f_reg[5][22]  ( .CLK(n5908), .D(N10340), .Q(
        decodedPacket5_o[22]) );
  LATCHX1 \decodedPacket_f_reg[5][21]  ( .CLK(n5908), .D(N10339), .Q(
        decodedPacket5_o[21]) );
  LATCHX1 \decodedPacket_f_reg[5][20]  ( .CLK(n5908), .D(N10338), .Q(
        decodedPacket5_o[20]) );
  LATCHX1 \decodedPacket_f_reg[5][19]  ( .CLK(n5908), .D(N10337), .Q(
        decodedPacket5_o[19]) );
  LATCHX1 \decodedPacket_f_reg[5][18]  ( .CLK(n5908), .D(N10336), .Q(
        decodedPacket5_o[18]) );
  LATCHX1 \decodedPacket_f_reg[5][17]  ( .CLK(n5908), .D(N10335), .Q(
        decodedPacket5_o[17]) );
  LATCHX1 \decodedPacket_f_reg[5][16]  ( .CLK(n5908), .D(N10334), .Q(
        decodedPacket5_o[16]) );
  LATCHX1 \decodedPacket_f_reg[5][15]  ( .CLK(n5908), .D(N10333), .Q(
        decodedPacket5_o[15]) );
  LATCHX1 \decodedPacket_f_reg[5][14]  ( .CLK(n5908), .D(N10332), .Q(
        decodedPacket5_o[14]) );
  LATCHX1 \decodedPacket_f_reg[5][13]  ( .CLK(n5908), .D(N10331), .Q(
        decodedPacket5_o[13]) );
  LATCHX1 \decodedPacket_f_reg[5][12]  ( .CLK(n5908), .D(N10330), .Q(
        decodedPacket5_o[12]) );
  LATCHX1 \decodedPacket_f_reg[5][11]  ( .CLK(n5907), .D(N10329), .Q(
        decodedPacket5_o[11]) );
  LATCHX1 \decodedPacket_f_reg[5][10]  ( .CLK(n5907), .D(N10328), .Q(
        decodedPacket5_o[10]) );
  LATCHX1 \decodedPacket_f_reg[5][9]  ( .CLK(n5907), .D(N10327), .Q(
        decodedPacket5_o[9]) );
  LATCHX1 \decodedPacket_f_reg[5][8]  ( .CLK(n5907), .D(N10326), .Q(
        decodedPacket5_o[8]) );
  LATCHX1 \decodedPacket_f_reg[5][7]  ( .CLK(n5907), .D(N10325), .Q(
        decodedPacket5_o[7]) );
  LATCHX1 \decodedPacket_f_reg[5][6]  ( .CLK(n5907), .D(N10324), .Q(
        decodedPacket5_o[6]) );
  LATCHX1 \decodedPacket_f_reg[5][5]  ( .CLK(n5907), .D(N10323), .Q(
        decodedPacket5_o[5]) );
  LATCHX1 \decodedPacket_f_reg[5][4]  ( .CLK(n5907), .D(N10322), .Q(
        decodedPacket5_o[4]) );
  LATCHX1 \decodedPacket_f_reg[5][3]  ( .CLK(n5907), .D(N10321), .Q(
        decodedPacket5_o[3]) );
  LATCHX1 \decodedPacket_f_reg[5][2]  ( .CLK(n5907), .D(N10320), .Q(
        decodedPacket5_o[2]) );
  LATCHX1 \decodedPacket_f_reg[5][1]  ( .CLK(n5907), .D(N10319), .Q(
        decodedPacket5_o[1]) );
  LATCHX1 \decodedPacket_f_reg[5][0]  ( .CLK(n5907), .D(N10318), .Q(
        decodedPacket5_o[0]) );
  LATCHX1 \decodedPacket_f_reg[4][121]  ( .CLK(n5901), .D(N10312), .Q(
        decodedPacket4_o[121]) );
  LATCHX1 \decodedPacket_f_reg[4][120]  ( .CLK(n5902), .D(N10311), .Q(
        decodedPacket4_o[120]) );
  LATCHX1 \decodedPacket_f_reg[4][119]  ( .CLK(n5906), .D(N10310), .Q(
        decodedPacket4_o[119]) );
  LATCHX1 \decodedPacket_f_reg[4][118]  ( .CLK(n5906), .D(N10309), .Q(
        decodedPacket4_o[118]) );
  LATCHX1 \decodedPacket_f_reg[4][117]  ( .CLK(n5906), .D(N10308), .Q(
        decodedPacket4_o[117]) );
  LATCHX1 \decodedPacket_f_reg[4][116]  ( .CLK(n5906), .D(N10307), .Q(
        decodedPacket4_o[116]) );
  LATCHX1 \decodedPacket_f_reg[4][115]  ( .CLK(n5906), .D(N10306), .Q(
        decodedPacket4_o[115]) );
  LATCHX1 \decodedPacket_f_reg[4][114]  ( .CLK(n5906), .D(N10305), .Q(
        decodedPacket4_o[114]) );
  LATCHX1 \decodedPacket_f_reg[4][113]  ( .CLK(n5906), .D(N10304), .Q(
        decodedPacket4_o[113]) );
  LATCHX1 \decodedPacket_f_reg[4][112]  ( .CLK(n5906), .D(N10303), .Q(
        decodedPacket4_o[112]) );
  LATCHX1 \decodedPacket_f_reg[4][111]  ( .CLK(n5906), .D(N10302), .Q(
        decodedPacket4_o[111]) );
  LATCHX1 \decodedPacket_f_reg[4][110]  ( .CLK(n5906), .D(N10301), .Q(
        decodedPacket4_o[110]) );
  LATCHX1 \decodedPacket_f_reg[4][109]  ( .CLK(n5906), .D(N10300), .Q(
        decodedPacket4_o[109]) );
  LATCHX1 \decodedPacket_f_reg[4][108]  ( .CLK(n5906), .D(N10299), .Q(
        decodedPacket4_o[108]) );
  LATCHX1 \decodedPacket_f_reg[4][107]  ( .CLK(n5905), .D(N10298), .Q(
        decodedPacket4_o[107]) );
  LATCHX1 \decodedPacket_f_reg[4][106]  ( .CLK(n5905), .D(N10297), .Q(
        decodedPacket4_o[106]) );
  LATCHX1 \decodedPacket_f_reg[4][105]  ( .CLK(n5905), .D(N10296), .Q(
        decodedPacket4_o[105]) );
  LATCHX1 \decodedPacket_f_reg[4][104]  ( .CLK(n5905), .D(N10295), .Q(
        decodedPacket4_o[104]) );
  LATCHX1 \decodedPacket_f_reg[4][103]  ( .CLK(n5905), .D(N10294), .Q(
        decodedPacket4_o[103]) );
  LATCHX1 \decodedPacket_f_reg[4][102]  ( .CLK(n5905), .D(N10293), .Q(
        decodedPacket4_o[102]) );
  LATCHX1 \decodedPacket_f_reg[4][101]  ( .CLK(n5905), .D(N10292), .Q(
        decodedPacket4_o[101]) );
  LATCHX1 \decodedPacket_f_reg[4][100]  ( .CLK(n5905), .D(N10291), .Q(
        decodedPacket4_o[100]) );
  LATCHX1 \decodedPacket_f_reg[4][99]  ( .CLK(n5905), .D(N10290), .Q(
        decodedPacket4_o[99]) );
  LATCHX1 \decodedPacket_f_reg[4][98]  ( .CLK(n5905), .D(N10288), .Q(
        decodedPacket4_o[98]) );
  LATCHX1 \decodedPacket_f_reg[4][97]  ( .CLK(n5905), .D(N10286), .Q(
        decodedPacket4_o[97]) );
  LATCHX1 \decodedPacket_f_reg[4][96]  ( .CLK(n5905), .D(N10285), .Q(
        decodedPacket4_o[96]) );
  LATCHX1 \decodedPacket_f_reg[4][95]  ( .CLK(n5904), .D(N10284), .Q(
        decodedPacket4_o[95]) );
  LATCHX1 \decodedPacket_f_reg[4][94]  ( .CLK(n5904), .D(N10283), .Q(
        decodedPacket4_o[94]) );
  LATCHX1 \decodedPacket_f_reg[4][93]  ( .CLK(n5904), .D(N10282), .Q(
        decodedPacket4_o[93]) );
  LATCHX1 \decodedPacket_f_reg[4][92]  ( .CLK(n5904), .D(N10281), .Q(
        decodedPacket4_o[92]) );
  LATCHX1 \decodedPacket_f_reg[4][91]  ( .CLK(n5904), .D(N10280), .Q(
        decodedPacket4_o[91]) );
  LATCHX1 \decodedPacket_f_reg[4][90]  ( .CLK(n5904), .D(N10279), .Q(
        decodedPacket4_o[90]) );
  LATCHX1 \decodedPacket_f_reg[4][89]  ( .CLK(n5904), .D(N10278), .Q(
        decodedPacket4_o[89]) );
  LATCHX1 \decodedPacket_f_reg[4][88]  ( .CLK(n5904), .D(N10277), .Q(
        decodedPacket4_o[88]) );
  LATCHX1 \decodedPacket_f_reg[4][87]  ( .CLK(n5904), .D(N10276), .Q(
        decodedPacket4_o[87]) );
  LATCHX1 \decodedPacket_f_reg[4][86]  ( .CLK(n5904), .D(N10275), .Q(
        decodedPacket4_o[86]) );
  LATCHX1 \decodedPacket_f_reg[4][85]  ( .CLK(n5904), .D(N10274), .Q(
        decodedPacket4_o[85]) );
  LATCHX1 \decodedPacket_f_reg[4][84]  ( .CLK(n5904), .D(N10273), .Q(
        decodedPacket4_o[84]) );
  LATCHX1 \decodedPacket_f_reg[4][83]  ( .CLK(n5903), .D(N10272), .Q(
        decodedPacket4_o[83]) );
  LATCHX1 \decodedPacket_f_reg[4][82]  ( .CLK(n5903), .D(N10271), .Q(
        decodedPacket4_o[82]) );
  LATCHX1 \decodedPacket_f_reg[4][81]  ( .CLK(n5903), .D(N10270), .Q(
        decodedPacket4_o[81]) );
  LATCHX1 \decodedPacket_f_reg[4][80]  ( .CLK(n5903), .D(N10269), .Q(
        decodedPacket4_o[80]) );
  LATCHX1 \decodedPacket_f_reg[4][79]  ( .CLK(n5903), .D(N10268), .Q(
        decodedPacket4_o[79]) );
  LATCHX1 \decodedPacket_f_reg[4][78]  ( .CLK(n5903), .D(N10267), .Q(
        decodedPacket4_o[78]) );
  LATCHX1 \decodedPacket_f_reg[4][77]  ( .CLK(n5903), .D(N10266), .Q(
        decodedPacket4_o[77]) );
  LATCHX1 \decodedPacket_f_reg[4][76]  ( .CLK(n5903), .D(N10265), .Q(
        decodedPacket4_o[76]) );
  LATCHX1 \decodedPacket_f_reg[4][75]  ( .CLK(n5903), .D(N10264), .Q(
        decodedPacket4_o[75]) );
  LATCHX1 \decodedPacket_f_reg[4][74]  ( .CLK(n5903), .D(N10263), .Q(
        decodedPacket4_o[74]) );
  LATCHX1 \decodedPacket_f_reg[4][73]  ( .CLK(n5903), .D(N10262), .Q(
        decodedPacket4_o[73]) );
  LATCHX1 \decodedPacket_f_reg[4][72]  ( .CLK(n5903), .D(N10261), .Q(
        decodedPacket4_o[72]) );
  LATCHX1 \decodedPacket_f_reg[4][71]  ( .CLK(n5902), .D(N10260), .Q(
        decodedPacket4_o[71]) );
  LATCHX1 \decodedPacket_f_reg[4][70]  ( .CLK(n5902), .D(N10259), .Q(
        decodedPacket4_o[70]) );
  LATCHX1 \decodedPacket_f_reg[4][69]  ( .CLK(n5902), .D(N10258), .Q(
        decodedPacket4_o[69]) );
  LATCHX1 \decodedPacket_f_reg[4][68]  ( .CLK(n5902), .D(N10257), .Q(
        decodedPacket4_o[68]) );
  LATCHX1 \decodedPacket_f_reg[4][67]  ( .CLK(n5902), .D(N10256), .Q(
        decodedPacket4_o[67]) );
  LATCHX1 \decodedPacket_f_reg[4][66]  ( .CLK(n5902), .D(N10255), .Q(
        decodedPacket4_o[66]) );
  LATCHX1 \decodedPacket_f_reg[4][65]  ( .CLK(n5902), .D(N10254), .Q(
        decodedPacket4_o[65]) );
  LATCHX1 \decodedPacket_f_reg[4][64]  ( .CLK(n5902), .D(N10253), .Q(
        decodedPacket4_o[64]) );
  LATCHX1 \decodedPacket_f_reg[4][63]  ( .CLK(n5902), .D(N10252), .Q(
        decodedPacket4_o[63]) );
  LATCHX1 \decodedPacket_f_reg[4][62]  ( .CLK(n5902), .D(N10251), .Q(
        decodedPacket4_o[62]) );
  LATCHX1 \decodedPacket_f_reg[4][61]  ( .CLK(n5902), .D(N10250), .Q(
        decodedPacket4_o[61]) );
  LATCHX1 \decodedPacket_f_reg[4][60]  ( .CLK(n5902), .D(N10249), .Q(
        decodedPacket4_o[60]) );
  LATCHX1 \decodedPacket_f_reg[4][59]  ( .CLK(n5901), .D(N10248), .Q(
        decodedPacket4_o[59]) );
  LATCHX1 \decodedPacket_f_reg[4][58]  ( .CLK(n5901), .D(N10247), .Q(
        decodedPacket4_o[58]) );
  LATCHX1 \decodedPacket_f_reg[4][57]  ( .CLK(n5901), .D(N10246), .Q(
        decodedPacket4_o[57]) );
  LATCHX1 \decodedPacket_f_reg[4][56]  ( .CLK(n5901), .D(N10245), .Q(
        decodedPacket4_o[56]) );
  LATCHX1 \decodedPacket_f_reg[4][55]  ( .CLK(n5901), .D(N10244), .Q(
        decodedPacket4_o[55]) );
  LATCHX1 \decodedPacket_f_reg[4][54]  ( .CLK(n5901), .D(N10243), .Q(
        decodedPacket4_o[54]) );
  LATCHX1 \decodedPacket_f_reg[4][53]  ( .CLK(n5901), .D(N10242), .Q(
        decodedPacket4_o[53]) );
  LATCHX1 \decodedPacket_f_reg[4][52]  ( .CLK(n5901), .D(N10241), .Q(
        decodedPacket4_o[52]) );
  LATCHX1 \decodedPacket_f_reg[4][51]  ( .CLK(n5901), .D(N10240), .Q(
        decodedPacket4_o[51]) );
  LATCHX1 \decodedPacket_f_reg[4][50]  ( .CLK(n5901), .D(N10239), .Q(
        decodedPacket4_o[50]) );
  LATCHX1 \decodedPacket_f_reg[4][49]  ( .CLK(n5901), .D(N10238), .Q(
        decodedPacket4_o[49]) );
  LATCHX1 \decodedPacket_f_reg[4][48]  ( .CLK(n5901), .D(N10236), .Q(
        decodedPacket4_o[48]) );
  LATCHX1 \decodedPacket_f_reg[4][47]  ( .CLK(n5900), .D(N10235), .Q(
        decodedPacket4_o[47]) );
  LATCHX1 \decodedPacket_f_reg[4][46]  ( .CLK(n5900), .D(N10234), .Q(
        decodedPacket4_o[46]) );
  LATCHX1 \decodedPacket_f_reg[4][45]  ( .CLK(n5900), .D(N10233), .Q(
        decodedPacket4_o[45]) );
  LATCHX1 \decodedPacket_f_reg[4][44]  ( .CLK(n5900), .D(N10232), .Q(
        decodedPacket4_o[44]) );
  LATCHX1 \decodedPacket_f_reg[4][43]  ( .CLK(n5900), .D(N10231), .Q(
        decodedPacket4_o[43]) );
  LATCHX1 \decodedPacket_f_reg[4][42]  ( .CLK(n5900), .D(N10230), .Q(
        decodedPacket4_o[42]) );
  LATCHX1 \decodedPacket_f_reg[4][41]  ( .CLK(n5900), .D(N10229), .Q(
        decodedPacket4_o[41]) );
  LATCHX1 \decodedPacket_f_reg[4][40]  ( .CLK(n5900), .D(N10228), .Q(
        decodedPacket4_o[40]) );
  LATCHX1 \decodedPacket_f_reg[4][39]  ( .CLK(n5900), .D(N10227), .Q(
        decodedPacket4_o[39]) );
  LATCHX1 \decodedPacket_f_reg[4][38]  ( .CLK(n5900), .D(N10226), .Q(
        decodedPacket4_o[38]) );
  LATCHX1 \decodedPacket_f_reg[4][37]  ( .CLK(n5900), .D(N10225), .Q(
        decodedPacket4_o[37]) );
  LATCHX1 \decodedPacket_f_reg[4][36]  ( .CLK(n5900), .D(N10224), .Q(
        decodedPacket4_o[36]) );
  LATCHX1 \decodedPacket_f_reg[4][35]  ( .CLK(n5899), .D(N10223), .Q(
        decodedPacket4_o[35]) );
  LATCHX1 \decodedPacket_f_reg[4][34]  ( .CLK(n5899), .D(N10222), .Q(
        decodedPacket4_o[34]) );
  LATCHX1 \decodedPacket_f_reg[4][33]  ( .CLK(n5899), .D(N10221), .Q(
        decodedPacket4_o[33]) );
  LATCHX1 \decodedPacket_f_reg[4][32]  ( .CLK(n5899), .D(N10220), .Q(
        decodedPacket4_o[32]) );
  LATCHX1 \decodedPacket_f_reg[4][31]  ( .CLK(n5899), .D(N10219), .Q(
        decodedPacket4_o[31]) );
  LATCHX1 \decodedPacket_f_reg[4][30]  ( .CLK(n5899), .D(N10218), .Q(
        decodedPacket4_o[30]) );
  LATCHX1 \decodedPacket_f_reg[4][29]  ( .CLK(n5899), .D(N10217), .Q(
        decodedPacket4_o[29]) );
  LATCHX1 \decodedPacket_f_reg[4][28]  ( .CLK(n5899), .D(N10216), .Q(
        decodedPacket4_o[28]) );
  LATCHX1 \decodedPacket_f_reg[4][27]  ( .CLK(n5899), .D(N10215), .Q(
        decodedPacket4_o[27]) );
  LATCHX1 \decodedPacket_f_reg[4][26]  ( .CLK(n5899), .D(N10214), .Q(
        decodedPacket4_o[26]) );
  LATCHX1 \decodedPacket_f_reg[4][25]  ( .CLK(n5899), .D(N10213), .Q(
        decodedPacket4_o[25]) );
  LATCHX1 \decodedPacket_f_reg[4][24]  ( .CLK(n5899), .D(N10212), .Q(
        decodedPacket4_o[24]) );
  LATCHX1 \decodedPacket_f_reg[4][23]  ( .CLK(n5898), .D(N10211), .Q(
        decodedPacket4_o[23]) );
  LATCHX1 \decodedPacket_f_reg[4][22]  ( .CLK(n5898), .D(N10210), .Q(
        decodedPacket4_o[22]) );
  LATCHX1 \decodedPacket_f_reg[4][21]  ( .CLK(n5898), .D(N10209), .Q(
        decodedPacket4_o[21]) );
  LATCHX1 \decodedPacket_f_reg[4][20]  ( .CLK(n5898), .D(N10208), .Q(
        decodedPacket4_o[20]) );
  LATCHX1 \decodedPacket_f_reg[4][19]  ( .CLK(n5898), .D(N10207), .Q(
        decodedPacket4_o[19]) );
  LATCHX1 \decodedPacket_f_reg[4][18]  ( .CLK(n5898), .D(N10206), .Q(
        decodedPacket4_o[18]) );
  LATCHX1 \decodedPacket_f_reg[4][17]  ( .CLK(n5898), .D(N10205), .Q(
        decodedPacket4_o[17]) );
  LATCHX1 \decodedPacket_f_reg[4][16]  ( .CLK(n5898), .D(N10204), .Q(
        decodedPacket4_o[16]) );
  LATCHX1 \decodedPacket_f_reg[4][15]  ( .CLK(n5898), .D(N10203), .Q(
        decodedPacket4_o[15]) );
  LATCHX1 \decodedPacket_f_reg[4][14]  ( .CLK(n5898), .D(N10202), .Q(
        decodedPacket4_o[14]) );
  LATCHX1 \decodedPacket_f_reg[4][13]  ( .CLK(n5898), .D(N10201), .Q(
        decodedPacket4_o[13]) );
  LATCHX1 \decodedPacket_f_reg[4][12]  ( .CLK(n5898), .D(N10200), .Q(
        decodedPacket4_o[12]) );
  LATCHX1 \decodedPacket_f_reg[4][11]  ( .CLK(n5897), .D(N10199), .Q(
        decodedPacket4_o[11]) );
  LATCHX1 \decodedPacket_f_reg[4][10]  ( .CLK(n5897), .D(N10198), .Q(
        decodedPacket4_o[10]) );
  LATCHX1 \decodedPacket_f_reg[4][9]  ( .CLK(n5897), .D(N10197), .Q(
        decodedPacket4_o[9]) );
  LATCHX1 \decodedPacket_f_reg[4][8]  ( .CLK(n5897), .D(N10196), .Q(
        decodedPacket4_o[8]) );
  LATCHX1 \decodedPacket_f_reg[4][7]  ( .CLK(n5897), .D(N10195), .Q(
        decodedPacket4_o[7]) );
  LATCHX1 \decodedPacket_f_reg[4][6]  ( .CLK(n5897), .D(N10194), .Q(
        decodedPacket4_o[6]) );
  LATCHX1 \decodedPacket_f_reg[4][5]  ( .CLK(n5897), .D(N10193), .Q(
        decodedPacket4_o[5]) );
  LATCHX1 \decodedPacket_f_reg[4][4]  ( .CLK(n5897), .D(N10192), .Q(
        decodedPacket4_o[4]) );
  LATCHX1 \decodedPacket_f_reg[4][3]  ( .CLK(n5897), .D(N10191), .Q(
        decodedPacket4_o[3]) );
  LATCHX1 \decodedPacket_f_reg[4][2]  ( .CLK(n5897), .D(N10190), .Q(
        decodedPacket4_o[2]) );
  LATCHX1 \decodedPacket_f_reg[4][1]  ( .CLK(n5897), .D(N10189), .Q(
        decodedPacket4_o[1]) );
  LATCHX1 \decodedPacket_f_reg[4][0]  ( .CLK(n5897), .D(N10188), .Q(
        decodedPacket4_o[0]) );
  LATCHX1 \decodedPacket_f_reg[3][121]  ( .CLK(n5891), .D(N10182), .Q(
        decodedPacket3_o[121]) );
  LATCHX1 \decodedPacket_f_reg[3][120]  ( .CLK(n5892), .D(N10181), .Q(
        decodedPacket3_o[120]) );
  LATCHX1 \decodedPacket_f_reg[3][119]  ( .CLK(n5896), .D(N10180), .Q(
        decodedPacket3_o[119]) );
  LATCHX1 \decodedPacket_f_reg[3][118]  ( .CLK(n5896), .D(N10179), .Q(
        decodedPacket3_o[118]) );
  LATCHX1 \decodedPacket_f_reg[3][117]  ( .CLK(n5896), .D(N10178), .Q(
        decodedPacket3_o[117]) );
  LATCHX1 \decodedPacket_f_reg[3][116]  ( .CLK(n5896), .D(N10177), .Q(
        decodedPacket3_o[116]) );
  LATCHX1 \decodedPacket_f_reg[3][115]  ( .CLK(n5896), .D(N10176), .Q(
        decodedPacket3_o[115]) );
  LATCHX1 \decodedPacket_f_reg[3][114]  ( .CLK(n5896), .D(N10175), .Q(
        decodedPacket3_o[114]) );
  LATCHX1 \decodedPacket_f_reg[3][113]  ( .CLK(n5896), .D(N10174), .Q(
        decodedPacket3_o[113]) );
  LATCHX1 \decodedPacket_f_reg[3][112]  ( .CLK(n5896), .D(N10173), .Q(
        decodedPacket3_o[112]) );
  LATCHX1 \decodedPacket_f_reg[3][111]  ( .CLK(n5896), .D(N10172), .Q(
        decodedPacket3_o[111]) );
  LATCHX1 \decodedPacket_f_reg[3][110]  ( .CLK(n5896), .D(N10171), .Q(
        decodedPacket3_o[110]) );
  LATCHX1 \decodedPacket_f_reg[3][109]  ( .CLK(n5896), .D(N10170), .Q(
        decodedPacket3_o[109]) );
  LATCHX1 \decodedPacket_f_reg[3][108]  ( .CLK(n5896), .D(N10169), .Q(
        decodedPacket3_o[108]) );
  LATCHX1 \decodedPacket_f_reg[3][107]  ( .CLK(n5895), .D(N10168), .Q(
        decodedPacket3_o[107]) );
  LATCHX1 \decodedPacket_f_reg[3][106]  ( .CLK(n5895), .D(N10167), .Q(
        decodedPacket3_o[106]) );
  LATCHX1 \decodedPacket_f_reg[3][105]  ( .CLK(n5895), .D(N10166), .Q(
        decodedPacket3_o[105]) );
  LATCHX1 \decodedPacket_f_reg[3][104]  ( .CLK(n5895), .D(N10165), .Q(
        decodedPacket3_o[104]) );
  LATCHX1 \decodedPacket_f_reg[3][103]  ( .CLK(n5895), .D(N10164), .Q(
        decodedPacket3_o[103]) );
  LATCHX1 \decodedPacket_f_reg[3][102]  ( .CLK(n5895), .D(N10163), .Q(
        decodedPacket3_o[102]) );
  LATCHX1 \decodedPacket_f_reg[3][101]  ( .CLK(n5895), .D(N10162), .Q(
        decodedPacket3_o[101]) );
  LATCHX1 \decodedPacket_f_reg[3][100]  ( .CLK(n5895), .D(N10161), .Q(
        decodedPacket3_o[100]) );
  LATCHX1 \decodedPacket_f_reg[3][99]  ( .CLK(n5895), .D(N10160), .Q(
        decodedPacket3_o[99]) );
  LATCHX1 \decodedPacket_f_reg[3][98]  ( .CLK(n5895), .D(N10158), .Q(
        decodedPacket3_o[98]) );
  LATCHX1 \decodedPacket_f_reg[3][97]  ( .CLK(n5895), .D(N10156), .Q(
        decodedPacket3_o[97]) );
  LATCHX1 \decodedPacket_f_reg[3][96]  ( .CLK(n5895), .D(N10155), .Q(
        decodedPacket3_o[96]) );
  LATCHX1 \decodedPacket_f_reg[3][95]  ( .CLK(n5894), .D(N10154), .Q(
        decodedPacket3_o[95]) );
  LATCHX1 \decodedPacket_f_reg[3][94]  ( .CLK(n5894), .D(N10153), .Q(
        decodedPacket3_o[94]) );
  LATCHX1 \decodedPacket_f_reg[3][93]  ( .CLK(n5894), .D(N10152), .Q(
        decodedPacket3_o[93]) );
  LATCHX1 \decodedPacket_f_reg[3][92]  ( .CLK(n5894), .D(N10151), .Q(
        decodedPacket3_o[92]) );
  LATCHX1 \decodedPacket_f_reg[3][91]  ( .CLK(n5894), .D(N10150), .Q(
        decodedPacket3_o[91]) );
  LATCHX1 \decodedPacket_f_reg[3][90]  ( .CLK(n5894), .D(N10149), .Q(
        decodedPacket3_o[90]) );
  LATCHX1 \decodedPacket_f_reg[3][89]  ( .CLK(n5894), .D(N10148), .Q(
        decodedPacket3_o[89]) );
  LATCHX1 \decodedPacket_f_reg[3][88]  ( .CLK(n5894), .D(N10147), .Q(
        decodedPacket3_o[88]) );
  LATCHX1 \decodedPacket_f_reg[3][87]  ( .CLK(n5894), .D(N10146), .Q(
        decodedPacket3_o[87]) );
  LATCHX1 \decodedPacket_f_reg[3][86]  ( .CLK(n5894), .D(N10145), .Q(
        decodedPacket3_o[86]) );
  LATCHX1 \decodedPacket_f_reg[3][85]  ( .CLK(n5894), .D(N10144), .Q(
        decodedPacket3_o[85]) );
  LATCHX1 \decodedPacket_f_reg[3][84]  ( .CLK(n5894), .D(N10143), .Q(
        decodedPacket3_o[84]) );
  LATCHX1 \decodedPacket_f_reg[3][83]  ( .CLK(n5893), .D(N10142), .Q(
        decodedPacket3_o[83]) );
  LATCHX1 \decodedPacket_f_reg[3][82]  ( .CLK(n5893), .D(N10141), .Q(
        decodedPacket3_o[82]) );
  LATCHX1 \decodedPacket_f_reg[3][81]  ( .CLK(n5893), .D(N10140), .Q(
        decodedPacket3_o[81]) );
  LATCHX1 \decodedPacket_f_reg[3][80]  ( .CLK(n5893), .D(N10139), .Q(
        decodedPacket3_o[80]) );
  LATCHX1 \decodedPacket_f_reg[3][79]  ( .CLK(n5893), .D(N10138), .Q(
        decodedPacket3_o[79]) );
  LATCHX1 \decodedPacket_f_reg[3][78]  ( .CLK(n5893), .D(N10137), .Q(
        decodedPacket3_o[78]) );
  LATCHX1 \decodedPacket_f_reg[3][77]  ( .CLK(n5893), .D(N10136), .Q(
        decodedPacket3_o[77]) );
  LATCHX1 \decodedPacket_f_reg[3][76]  ( .CLK(n5893), .D(N10135), .Q(
        decodedPacket3_o[76]) );
  LATCHX1 \decodedPacket_f_reg[3][75]  ( .CLK(n5893), .D(N10134), .Q(
        decodedPacket3_o[75]) );
  LATCHX1 \decodedPacket_f_reg[3][74]  ( .CLK(n5893), .D(N10133), .Q(
        decodedPacket3_o[74]) );
  LATCHX1 \decodedPacket_f_reg[3][73]  ( .CLK(n5893), .D(N10132), .Q(
        decodedPacket3_o[73]) );
  LATCHX1 \decodedPacket_f_reg[3][72]  ( .CLK(n5893), .D(N10131), .Q(
        decodedPacket3_o[72]) );
  LATCHX1 \decodedPacket_f_reg[3][71]  ( .CLK(n5892), .D(N10130), .Q(
        decodedPacket3_o[71]) );
  LATCHX1 \decodedPacket_f_reg[3][70]  ( .CLK(n5892), .D(N10129), .Q(
        decodedPacket3_o[70]) );
  LATCHX1 \decodedPacket_f_reg[3][69]  ( .CLK(n5892), .D(N10128), .Q(
        decodedPacket3_o[69]) );
  LATCHX1 \decodedPacket_f_reg[3][68]  ( .CLK(n5892), .D(N10127), .Q(
        decodedPacket3_o[68]) );
  LATCHX1 \decodedPacket_f_reg[3][67]  ( .CLK(n5892), .D(N10126), .Q(
        decodedPacket3_o[67]) );
  LATCHX1 \decodedPacket_f_reg[3][66]  ( .CLK(n5892), .D(N10125), .Q(
        decodedPacket3_o[66]) );
  LATCHX1 \decodedPacket_f_reg[3][65]  ( .CLK(n5892), .D(N10124), .Q(
        decodedPacket3_o[65]) );
  LATCHX1 \decodedPacket_f_reg[3][64]  ( .CLK(n5892), .D(N10123), .Q(
        decodedPacket3_o[64]) );
  LATCHX1 \decodedPacket_f_reg[3][63]  ( .CLK(n5892), .D(N10122), .Q(
        decodedPacket3_o[63]) );
  LATCHX1 \decodedPacket_f_reg[3][62]  ( .CLK(n5892), .D(N10121), .Q(
        decodedPacket3_o[62]) );
  LATCHX1 \decodedPacket_f_reg[3][61]  ( .CLK(n5892), .D(N10120), .Q(
        decodedPacket3_o[61]) );
  LATCHX1 \decodedPacket_f_reg[3][60]  ( .CLK(n5892), .D(N10119), .Q(
        decodedPacket3_o[60]) );
  LATCHX1 \decodedPacket_f_reg[3][59]  ( .CLK(n5891), .D(N10118), .Q(
        decodedPacket3_o[59]) );
  LATCHX1 \decodedPacket_f_reg[3][58]  ( .CLK(n5891), .D(N10117), .Q(
        decodedPacket3_o[58]) );
  LATCHX1 \decodedPacket_f_reg[3][57]  ( .CLK(n5891), .D(N10116), .Q(
        decodedPacket3_o[57]) );
  LATCHX1 \decodedPacket_f_reg[3][56]  ( .CLK(n5891), .D(N10115), .Q(
        decodedPacket3_o[56]) );
  LATCHX1 \decodedPacket_f_reg[3][55]  ( .CLK(n5891), .D(N10114), .Q(
        decodedPacket3_o[55]) );
  LATCHX1 \decodedPacket_f_reg[3][54]  ( .CLK(n5891), .D(N10113), .Q(
        decodedPacket3_o[54]) );
  LATCHX1 \decodedPacket_f_reg[3][53]  ( .CLK(n5891), .D(N10112), .Q(
        decodedPacket3_o[53]) );
  LATCHX1 \decodedPacket_f_reg[3][52]  ( .CLK(n5891), .D(N10111), .Q(
        decodedPacket3_o[52]) );
  LATCHX1 \decodedPacket_f_reg[3][51]  ( .CLK(n5891), .D(N10110), .Q(
        decodedPacket3_o[51]) );
  LATCHX1 \decodedPacket_f_reg[3][50]  ( .CLK(n5891), .D(N10109), .Q(
        decodedPacket3_o[50]) );
  LATCHX1 \decodedPacket_f_reg[3][49]  ( .CLK(n5891), .D(N10108), .Q(
        decodedPacket3_o[49]) );
  LATCHX1 \decodedPacket_f_reg[3][48]  ( .CLK(n5891), .D(N10106), .Q(
        decodedPacket3_o[48]) );
  LATCHX1 \decodedPacket_f_reg[3][47]  ( .CLK(n5890), .D(N10105), .Q(
        decodedPacket3_o[47]) );
  LATCHX1 \decodedPacket_f_reg[3][46]  ( .CLK(n5890), .D(N10104), .Q(
        decodedPacket3_o[46]) );
  LATCHX1 \decodedPacket_f_reg[3][45]  ( .CLK(n5890), .D(N10103), .Q(
        decodedPacket3_o[45]) );
  LATCHX1 \decodedPacket_f_reg[3][44]  ( .CLK(n5890), .D(N10102), .Q(
        decodedPacket3_o[44]) );
  LATCHX1 \decodedPacket_f_reg[3][43]  ( .CLK(n5890), .D(N10101), .Q(
        decodedPacket3_o[43]) );
  LATCHX1 \decodedPacket_f_reg[3][42]  ( .CLK(n5890), .D(N10100), .Q(
        decodedPacket3_o[42]) );
  LATCHX1 \decodedPacket_f_reg[3][41]  ( .CLK(n5890), .D(N10099), .Q(
        decodedPacket3_o[41]) );
  LATCHX1 \decodedPacket_f_reg[3][40]  ( .CLK(n5890), .D(N10098), .Q(
        decodedPacket3_o[40]) );
  LATCHX1 \decodedPacket_f_reg[3][39]  ( .CLK(n5890), .D(N10097), .Q(
        decodedPacket3_o[39]) );
  LATCHX1 \decodedPacket_f_reg[3][38]  ( .CLK(n5890), .D(N10096), .Q(
        decodedPacket3_o[38]) );
  LATCHX1 \decodedPacket_f_reg[3][37]  ( .CLK(n5890), .D(N10095), .Q(
        decodedPacket3_o[37]) );
  LATCHX1 \decodedPacket_f_reg[3][36]  ( .CLK(n5890), .D(N10094), .Q(
        decodedPacket3_o[36]) );
  LATCHX1 \decodedPacket_f_reg[3][35]  ( .CLK(n5889), .D(N10093), .Q(
        decodedPacket3_o[35]) );
  LATCHX1 \decodedPacket_f_reg[3][34]  ( .CLK(n5889), .D(N10092), .Q(
        decodedPacket3_o[34]) );
  LATCHX1 \decodedPacket_f_reg[3][33]  ( .CLK(n5889), .D(N10091), .Q(
        decodedPacket3_o[33]) );
  LATCHX1 \decodedPacket_f_reg[3][32]  ( .CLK(n5889), .D(N10090), .Q(
        decodedPacket3_o[32]) );
  LATCHX1 \decodedPacket_f_reg[3][31]  ( .CLK(n5889), .D(N10089), .Q(
        decodedPacket3_o[31]) );
  LATCHX1 \decodedPacket_f_reg[3][30]  ( .CLK(n5889), .D(N10088), .Q(
        decodedPacket3_o[30]) );
  LATCHX1 \decodedPacket_f_reg[3][29]  ( .CLK(n5889), .D(N10087), .Q(
        decodedPacket3_o[29]) );
  LATCHX1 \decodedPacket_f_reg[3][28]  ( .CLK(n5889), .D(N10086), .Q(
        decodedPacket3_o[28]) );
  LATCHX1 \decodedPacket_f_reg[3][27]  ( .CLK(n5889), .D(N10085), .Q(
        decodedPacket3_o[27]) );
  LATCHX1 \decodedPacket_f_reg[3][26]  ( .CLK(n5889), .D(N10084), .Q(
        decodedPacket3_o[26]) );
  LATCHX1 \decodedPacket_f_reg[3][25]  ( .CLK(n5889), .D(N10083), .Q(
        decodedPacket3_o[25]) );
  LATCHX1 \decodedPacket_f_reg[3][24]  ( .CLK(n5889), .D(N10082), .Q(
        decodedPacket3_o[24]) );
  LATCHX1 \decodedPacket_f_reg[3][23]  ( .CLK(n5888), .D(N10081), .Q(
        decodedPacket3_o[23]) );
  LATCHX1 \decodedPacket_f_reg[3][22]  ( .CLK(n5888), .D(N10080), .Q(
        decodedPacket3_o[22]) );
  LATCHX1 \decodedPacket_f_reg[3][21]  ( .CLK(n5888), .D(N10079), .Q(
        decodedPacket3_o[21]) );
  LATCHX1 \decodedPacket_f_reg[3][20]  ( .CLK(n5888), .D(N10078), .Q(
        decodedPacket3_o[20]) );
  LATCHX1 \decodedPacket_f_reg[3][19]  ( .CLK(n5888), .D(N10077), .Q(
        decodedPacket3_o[19]) );
  LATCHX1 \decodedPacket_f_reg[3][18]  ( .CLK(n5888), .D(N10076), .Q(
        decodedPacket3_o[18]) );
  LATCHX1 \decodedPacket_f_reg[3][17]  ( .CLK(n5888), .D(N10075), .Q(
        decodedPacket3_o[17]) );
  LATCHX1 \decodedPacket_f_reg[3][16]  ( .CLK(n5888), .D(N10074), .Q(
        decodedPacket3_o[16]) );
  LATCHX1 \decodedPacket_f_reg[3][15]  ( .CLK(n5888), .D(N10073), .Q(
        decodedPacket3_o[15]) );
  LATCHX1 \decodedPacket_f_reg[3][14]  ( .CLK(n5888), .D(N10072), .Q(
        decodedPacket3_o[14]) );
  LATCHX1 \decodedPacket_f_reg[3][13]  ( .CLK(n5888), .D(N10071), .Q(
        decodedPacket3_o[13]) );
  LATCHX1 \decodedPacket_f_reg[3][12]  ( .CLK(n5888), .D(N10070), .Q(
        decodedPacket3_o[12]) );
  LATCHX1 \decodedPacket_f_reg[3][11]  ( .CLK(n5887), .D(N10069), .Q(
        decodedPacket3_o[11]) );
  LATCHX1 \decodedPacket_f_reg[3][10]  ( .CLK(n5887), .D(N10068), .Q(
        decodedPacket3_o[10]) );
  LATCHX1 \decodedPacket_f_reg[3][9]  ( .CLK(n5887), .D(N10067), .Q(
        decodedPacket3_o[9]) );
  LATCHX1 \decodedPacket_f_reg[3][8]  ( .CLK(n5887), .D(N10066), .Q(
        decodedPacket3_o[8]) );
  LATCHX1 \decodedPacket_f_reg[3][7]  ( .CLK(n5887), .D(N10065), .Q(
        decodedPacket3_o[7]) );
  LATCHX1 \decodedPacket_f_reg[3][6]  ( .CLK(n5887), .D(N10064), .Q(
        decodedPacket3_o[6]) );
  LATCHX1 \decodedPacket_f_reg[3][5]  ( .CLK(n5887), .D(N10063), .Q(
        decodedPacket3_o[5]) );
  LATCHX1 \decodedPacket_f_reg[3][4]  ( .CLK(n5887), .D(N10062), .Q(
        decodedPacket3_o[4]) );
  LATCHX1 \decodedPacket_f_reg[3][3]  ( .CLK(n5887), .D(N10061), .Q(
        decodedPacket3_o[3]) );
  LATCHX1 \decodedPacket_f_reg[3][2]  ( .CLK(n5887), .D(N10060), .Q(
        decodedPacket3_o[2]) );
  LATCHX1 \decodedPacket_f_reg[3][1]  ( .CLK(n5887), .D(N10059), .Q(
        decodedPacket3_o[1]) );
  LATCHX1 \decodedPacket_f_reg[3][0]  ( .CLK(n5887), .D(N10058), .Q(
        decodedPacket3_o[0]) );
  LATCHX1 \decodedPacket_f_reg[2][121]  ( .CLK(n5877), .D(N10052), .Q(
        decodedPacket2_o[121]) );
  LATCHX1 \decodedPacket_f_reg[2][120]  ( .CLK(n5878), .D(N10051), .Q(
        decodedPacket2_o[120]) );
  LATCHX1 \decodedPacket_f_reg[2][119]  ( .CLK(n5886), .D(N10050), .Q(
        decodedPacket2_o[119]) );
  LATCHX1 \decodedPacket_f_reg[2][118]  ( .CLK(n5886), .D(N10049), .Q(
        decodedPacket2_o[118]) );
  LATCHX1 \decodedPacket_f_reg[2][117]  ( .CLK(n5886), .D(N10048), .Q(
        decodedPacket2_o[117]) );
  LATCHX1 \decodedPacket_f_reg[2][116]  ( .CLK(n5886), .D(N10047), .Q(
        decodedPacket2_o[116]) );
  LATCHX1 \decodedPacket_f_reg[2][115]  ( .CLK(n5886), .D(N10046), .Q(
        decodedPacket2_o[115]) );
  LATCHX1 \decodedPacket_f_reg[2][114]  ( .CLK(n5886), .D(N10045), .Q(
        decodedPacket2_o[114]) );
  LATCHX1 \decodedPacket_f_reg[2][113]  ( .CLK(n5886), .D(N10044), .Q(
        decodedPacket2_o[113]) );
  LATCHX1 \decodedPacket_f_reg[2][112]  ( .CLK(n5886), .D(N10043), .Q(
        decodedPacket2_o[112]) );
  LATCHX1 \decodedPacket_f_reg[2][111]  ( .CLK(n5886), .D(N10042), .Q(
        decodedPacket2_o[111]) );
  LATCHX1 \decodedPacket_f_reg[2][110]  ( .CLK(n5886), .D(N10041), .Q(
        decodedPacket2_o[110]) );
  LATCHX1 \decodedPacket_f_reg[2][109]  ( .CLK(n5886), .D(N10040), .Q(
        decodedPacket2_o[109]) );
  LATCHX1 \decodedPacket_f_reg[2][108]  ( .CLK(n5886), .D(N10039), .Q(
        decodedPacket2_o[108]) );
  LATCHX1 \decodedPacket_f_reg[2][107]  ( .CLK(n5885), .D(N10038), .Q(
        decodedPacket2_o[107]) );
  LATCHX1 \decodedPacket_f_reg[2][106]  ( .CLK(n5885), .D(N10037), .Q(
        decodedPacket2_o[106]) );
  LATCHX1 \decodedPacket_f_reg[2][105]  ( .CLK(n5885), .D(N10036), .Q(
        decodedPacket2_o[105]) );
  LATCHX1 \decodedPacket_f_reg[2][104]  ( .CLK(n5885), .D(N10035), .Q(
        decodedPacket2_o[104]) );
  LATCHX1 \decodedPacket_f_reg[2][103]  ( .CLK(n5885), .D(N10034), .Q(
        decodedPacket2_o[103]) );
  LATCHX1 \decodedPacket_f_reg[2][102]  ( .CLK(n5885), .D(N10033), .Q(
        decodedPacket2_o[102]) );
  LATCHX1 \decodedPacket_f_reg[2][101]  ( .CLK(n5885), .D(N10032), .Q(
        decodedPacket2_o[101]) );
  LATCHX1 \decodedPacket_f_reg[2][100]  ( .CLK(n5885), .D(N10031), .Q(
        decodedPacket2_o[100]) );
  LATCHX1 \decodedPacket_f_reg[2][99]  ( .CLK(n5885), .D(N10030), .Q(
        decodedPacket2_o[99]) );
  LATCHX1 \decodedPacket_f_reg[2][98]  ( .CLK(n5885), .D(N10028), .Q(
        decodedPacket2_o[98]) );
  LATCHX1 \decodedPacket_f_reg[2][97]  ( .CLK(n5885), .D(N10026), .Q(
        decodedPacket2_o[97]) );
  LATCHX1 \decodedPacket_f_reg[2][96]  ( .CLK(n5885), .D(N10025), .Q(
        decodedPacket2_o[96]) );
  LATCHX1 \decodedPacket_f_reg[2][95]  ( .CLK(n5884), .D(N10024), .Q(
        decodedPacket2_o[95]) );
  LATCHX1 \decodedPacket_f_reg[2][94]  ( .CLK(n5884), .D(N10023), .Q(
        decodedPacket2_o[94]) );
  LATCHX1 \decodedPacket_f_reg[2][93]  ( .CLK(n5884), .D(N10022), .Q(
        decodedPacket2_o[93]) );
  LATCHX1 \decodedPacket_f_reg[2][92]  ( .CLK(n5884), .D(N10021), .Q(
        decodedPacket2_o[92]) );
  LATCHX1 \decodedPacket_f_reg[2][91]  ( .CLK(n5884), .D(N10020), .Q(
        decodedPacket2_o[91]) );
  LATCHX1 \decodedPacket_f_reg[2][90]  ( .CLK(n5884), .D(N10019), .Q(
        decodedPacket2_o[90]) );
  LATCHX1 \decodedPacket_f_reg[2][89]  ( .CLK(n5884), .D(N10018), .Q(
        decodedPacket2_o[89]) );
  LATCHX1 \decodedPacket_f_reg[2][88]  ( .CLK(n5884), .D(N10017), .Q(
        decodedPacket2_o[88]) );
  LATCHX1 \decodedPacket_f_reg[2][87]  ( .CLK(n5884), .D(N10016), .Q(
        decodedPacket2_o[87]) );
  LATCHX1 \decodedPacket_f_reg[2][86]  ( .CLK(n5884), .D(N10015), .Q(
        decodedPacket2_o[86]) );
  LATCHX1 \decodedPacket_f_reg[2][85]  ( .CLK(n5884), .D(N10014), .Q(
        decodedPacket2_o[85]) );
  LATCHX1 \decodedPacket_f_reg[2][84]  ( .CLK(n5884), .D(N10013), .Q(
        decodedPacket2_o[84]) );
  LATCHX1 \decodedPacket_f_reg[2][83]  ( .CLK(n5883), .D(N10012), .Q(
        decodedPacket2_o[83]) );
  LATCHX1 \decodedPacket_f_reg[2][82]  ( .CLK(n5883), .D(N10011), .Q(
        decodedPacket2_o[82]) );
  LATCHX1 \decodedPacket_f_reg[2][81]  ( .CLK(n5883), .D(N10010), .Q(
        decodedPacket2_o[81]) );
  LATCHX1 \decodedPacket_f_reg[2][80]  ( .CLK(n5883), .D(N10009), .Q(
        decodedPacket2_o[80]) );
  LATCHX1 \decodedPacket_f_reg[2][79]  ( .CLK(n5883), .D(N10008), .Q(
        decodedPacket2_o[79]) );
  LATCHX1 \decodedPacket_f_reg[2][78]  ( .CLK(n5883), .D(N10007), .Q(
        decodedPacket2_o[78]) );
  LATCHX1 \decodedPacket_f_reg[2][77]  ( .CLK(n5883), .D(N10006), .Q(
        decodedPacket2_o[77]) );
  LATCHX1 \decodedPacket_f_reg[2][76]  ( .CLK(n5883), .D(N10005), .Q(
        decodedPacket2_o[76]) );
  LATCHX1 \decodedPacket_f_reg[2][75]  ( .CLK(n5883), .D(N10004), .Q(
        decodedPacket2_o[75]) );
  LATCHX1 \decodedPacket_f_reg[2][74]  ( .CLK(n5883), .D(N10003), .Q(
        decodedPacket2_o[74]) );
  LATCHX1 \decodedPacket_f_reg[2][73]  ( .CLK(n5883), .D(N10002), .Q(
        decodedPacket2_o[73]) );
  LATCHX1 \decodedPacket_f_reg[2][72]  ( .CLK(n5883), .D(N10001), .Q(
        decodedPacket2_o[72]) );
  LATCHX1 \decodedPacket_f_reg[2][71]  ( .CLK(n5882), .D(N10000), .Q(
        decodedPacket2_o[71]) );
  LATCHX1 \decodedPacket_f_reg[2][70]  ( .CLK(n5882), .D(N9999), .Q(
        decodedPacket2_o[70]) );
  LATCHX1 \decodedPacket_f_reg[2][69]  ( .CLK(n5882), .D(N9998), .Q(
        decodedPacket2_o[69]) );
  LATCHX1 \decodedPacket_f_reg[2][68]  ( .CLK(n5882), .D(N9997), .Q(
        decodedPacket2_o[68]) );
  LATCHX1 \decodedPacket_f_reg[2][67]  ( .CLK(n5882), .D(N9996), .Q(
        decodedPacket2_o[67]) );
  LATCHX1 \decodedPacket_f_reg[2][66]  ( .CLK(n5882), .D(N9995), .Q(
        decodedPacket2_o[66]) );
  LATCHX1 \decodedPacket_f_reg[2][65]  ( .CLK(n5882), .D(N9994), .Q(
        decodedPacket2_o[65]) );
  LATCHX1 \decodedPacket_f_reg[2][64]  ( .CLK(n5882), .D(N9993), .Q(
        decodedPacket2_o[64]) );
  LATCHX1 \decodedPacket_f_reg[2][63]  ( .CLK(n5882), .D(N9992), .Q(
        decodedPacket2_o[63]) );
  LATCHX1 \decodedPacket_f_reg[2][62]  ( .CLK(n5882), .D(N9991), .Q(
        decodedPacket2_o[62]) );
  LATCHX1 \decodedPacket_f_reg[2][61]  ( .CLK(n5882), .D(N9990), .Q(
        decodedPacket2_o[61]) );
  LATCHX1 \decodedPacket_f_reg[2][60]  ( .CLK(n5882), .D(N9989), .Q(
        decodedPacket2_o[60]) );
  LATCHX1 \decodedPacket_f_reg[2][59]  ( .CLK(n5881), .D(N9988), .Q(
        decodedPacket2_o[59]) );
  LATCHX1 \decodedPacket_f_reg[2][58]  ( .CLK(n5881), .D(N9987), .Q(
        decodedPacket2_o[58]) );
  LATCHX1 \decodedPacket_f_reg[2][57]  ( .CLK(n5881), .D(N9986), .Q(
        decodedPacket2_o[57]) );
  LATCHX1 \decodedPacket_f_reg[2][56]  ( .CLK(n5881), .D(N9985), .Q(
        decodedPacket2_o[56]) );
  LATCHX1 \decodedPacket_f_reg[2][55]  ( .CLK(n5881), .D(N9984), .Q(
        decodedPacket2_o[55]) );
  LATCHX1 \decodedPacket_f_reg[2][54]  ( .CLK(n5881), .D(N9983), .Q(
        decodedPacket2_o[54]) );
  LATCHX1 \decodedPacket_f_reg[2][53]  ( .CLK(n5881), .D(N9982), .Q(
        decodedPacket2_o[53]) );
  LATCHX1 \decodedPacket_f_reg[2][52]  ( .CLK(n5881), .D(N9981), .Q(
        decodedPacket2_o[52]) );
  LATCHX1 \decodedPacket_f_reg[2][51]  ( .CLK(n5881), .D(N9980), .Q(
        decodedPacket2_o[51]) );
  LATCHX1 \decodedPacket_f_reg[2][50]  ( .CLK(n5881), .D(N9979), .Q(
        decodedPacket2_o[50]) );
  LATCHX1 \decodedPacket_f_reg[2][49]  ( .CLK(n5881), .D(N9978), .Q(
        decodedPacket2_o[49]) );
  LATCHX1 \decodedPacket_f_reg[2][48]  ( .CLK(n5881), .D(N9976), .Q(
        decodedPacket2_o[48]) );
  LATCHX1 \decodedPacket_f_reg[2][47]  ( .CLK(n5880), .D(N9975), .Q(
        decodedPacket2_o[47]) );
  LATCHX1 \decodedPacket_f_reg[2][46]  ( .CLK(n5880), .D(N9974), .Q(
        decodedPacket2_o[46]) );
  LATCHX1 \decodedPacket_f_reg[2][45]  ( .CLK(n5880), .D(N9973), .Q(
        decodedPacket2_o[45]) );
  LATCHX1 \decodedPacket_f_reg[2][44]  ( .CLK(n5880), .D(N9972), .Q(
        decodedPacket2_o[44]) );
  LATCHX1 \decodedPacket_f_reg[2][43]  ( .CLK(n5880), .D(N9971), .Q(
        decodedPacket2_o[43]) );
  LATCHX1 \decodedPacket_f_reg[2][42]  ( .CLK(n5880), .D(N9970), .Q(
        decodedPacket2_o[42]) );
  LATCHX1 \decodedPacket_f_reg[2][41]  ( .CLK(n5880), .D(N9969), .Q(
        decodedPacket2_o[41]) );
  LATCHX1 \decodedPacket_f_reg[2][40]  ( .CLK(n5880), .D(N9968), .Q(
        decodedPacket2_o[40]) );
  LATCHX1 \decodedPacket_f_reg[2][39]  ( .CLK(n5880), .D(N9967), .Q(
        decodedPacket2_o[39]) );
  LATCHX1 \decodedPacket_f_reg[2][38]  ( .CLK(n5880), .D(N9966), .Q(
        decodedPacket2_o[38]) );
  LATCHX1 \decodedPacket_f_reg[2][37]  ( .CLK(n5880), .D(N9965), .Q(
        decodedPacket2_o[37]) );
  LATCHX1 \decodedPacket_f_reg[2][36]  ( .CLK(n5880), .D(N9964), .Q(
        decodedPacket2_o[36]) );
  LATCHX1 \decodedPacket_f_reg[2][35]  ( .CLK(n5879), .D(N9963), .Q(
        decodedPacket2_o[35]) );
  LATCHX1 \decodedPacket_f_reg[2][34]  ( .CLK(n5879), .D(N9962), .Q(
        decodedPacket2_o[34]) );
  LATCHX1 \decodedPacket_f_reg[2][33]  ( .CLK(n5879), .D(N9961), .Q(
        decodedPacket2_o[33]) );
  LATCHX1 \decodedPacket_f_reg[2][32]  ( .CLK(n5879), .D(N9960), .Q(
        decodedPacket2_o[32]) );
  LATCHX1 \decodedPacket_f_reg[2][31]  ( .CLK(n5879), .D(N9959), .Q(
        decodedPacket2_o[31]) );
  LATCHX1 \decodedPacket_f_reg[2][30]  ( .CLK(n5879), .D(N9958), .Q(
        decodedPacket2_o[30]) );
  LATCHX1 \decodedPacket_f_reg[2][29]  ( .CLK(n5879), .D(N9957), .Q(
        decodedPacket2_o[29]) );
  LATCHX1 \decodedPacket_f_reg[2][28]  ( .CLK(n5879), .D(N9956), .Q(
        decodedPacket2_o[28]) );
  LATCHX1 \decodedPacket_f_reg[2][27]  ( .CLK(n5879), .D(N9955), .Q(
        decodedPacket2_o[27]) );
  LATCHX1 \decodedPacket_f_reg[2][26]  ( .CLK(n5879), .D(N9954), .Q(
        decodedPacket2_o[26]) );
  LATCHX1 \decodedPacket_f_reg[2][25]  ( .CLK(n5879), .D(N9953), .Q(
        decodedPacket2_o[25]) );
  LATCHX1 \decodedPacket_f_reg[2][24]  ( .CLK(n5879), .D(N9952), .Q(
        decodedPacket2_o[24]) );
  LATCHX1 \decodedPacket_f_reg[2][23]  ( .CLK(n5878), .D(N9951), .Q(
        decodedPacket2_o[23]) );
  LATCHX1 \decodedPacket_f_reg[2][22]  ( .CLK(n5878), .D(N9950), .Q(
        decodedPacket2_o[22]) );
  LATCHX1 \decodedPacket_f_reg[2][21]  ( .CLK(n5878), .D(N9949), .Q(
        decodedPacket2_o[21]) );
  LATCHX1 \decodedPacket_f_reg[2][20]  ( .CLK(n5878), .D(N9948), .Q(
        decodedPacket2_o[20]) );
  LATCHX1 \decodedPacket_f_reg[2][19]  ( .CLK(n5878), .D(N9947), .Q(
        decodedPacket2_o[19]) );
  LATCHX1 \decodedPacket_f_reg[2][18]  ( .CLK(n5878), .D(N9946), .Q(
        decodedPacket2_o[18]) );
  LATCHX1 \decodedPacket_f_reg[2][17]  ( .CLK(n5878), .D(N9945), .Q(
        decodedPacket2_o[17]) );
  LATCHX1 \decodedPacket_f_reg[2][16]  ( .CLK(n5878), .D(N9944), .Q(
        decodedPacket2_o[16]) );
  LATCHX1 \decodedPacket_f_reg[2][15]  ( .CLK(n5878), .D(N9943), .Q(
        decodedPacket2_o[15]) );
  LATCHX1 \decodedPacket_f_reg[2][14]  ( .CLK(n5878), .D(N9942), .Q(
        decodedPacket2_o[14]) );
  LATCHX1 \decodedPacket_f_reg[2][13]  ( .CLK(n5878), .D(N9941), .Q(
        decodedPacket2_o[13]) );
  LATCHX1 \decodedPacket_f_reg[2][12]  ( .CLK(n5878), .D(N9940), .Q(
        decodedPacket2_o[12]) );
  LATCHX1 \decodedPacket_f_reg[2][11]  ( .CLK(n5877), .D(N9939), .Q(
        decodedPacket2_o[11]) );
  LATCHX1 \decodedPacket_f_reg[2][10]  ( .CLK(n5877), .D(N9938), .Q(
        decodedPacket2_o[10]) );
  LATCHX1 \decodedPacket_f_reg[2][9]  ( .CLK(n5877), .D(N9937), .Q(
        decodedPacket2_o[9]) );
  LATCHX1 \decodedPacket_f_reg[2][8]  ( .CLK(n5877), .D(N9936), .Q(
        decodedPacket2_o[8]) );
  LATCHX1 \decodedPacket_f_reg[2][7]  ( .CLK(n5877), .D(N9935), .Q(
        decodedPacket2_o[7]) );
  LATCHX1 \decodedPacket_f_reg[2][6]  ( .CLK(n5877), .D(N9934), .Q(
        decodedPacket2_o[6]) );
  LATCHX1 \decodedPacket_f_reg[2][5]  ( .CLK(n5877), .D(N9933), .Q(
        decodedPacket2_o[5]) );
  LATCHX1 \decodedPacket_f_reg[2][4]  ( .CLK(n5877), .D(N9932), .Q(
        decodedPacket2_o[4]) );
  LATCHX1 \decodedPacket_f_reg[2][3]  ( .CLK(n5877), .D(N9931), .Q(
        decodedPacket2_o[3]) );
  LATCHX1 \decodedPacket_f_reg[2][2]  ( .CLK(n5877), .D(N9930), .Q(
        decodedPacket2_o[2]) );
  LATCHX1 \decodedPacket_f_reg[2][1]  ( .CLK(n5877), .D(N9929), .Q(
        decodedPacket2_o[1]) );
  LATCHX1 \decodedPacket_f_reg[2][0]  ( .CLK(n5877), .D(N9928), .Q(
        decodedPacket2_o[0]) );
  LATCHX1 \decodedPacket_f_reg[1][121]  ( .CLK(n5871), .D(N9922), .Q(
        decodedPacket1_o[121]) );
  LATCHX1 \decodedPacket_f_reg[1][120]  ( .CLK(n5872), .D(N9921), .Q(
        decodedPacket1_o[120]) );
  LATCHX1 \decodedPacket_f_reg[1][119]  ( .CLK(n5876), .D(N9920), .Q(
        decodedPacket1_o[119]) );
  LATCHX1 \decodedPacket_f_reg[1][118]  ( .CLK(n5876), .D(N9919), .Q(
        decodedPacket1_o[118]) );
  LATCHX1 \decodedPacket_f_reg[1][117]  ( .CLK(n5876), .D(N9918), .Q(
        decodedPacket1_o[117]) );
  LATCHX1 \decodedPacket_f_reg[1][116]  ( .CLK(n5876), .D(N9917), .Q(
        decodedPacket1_o[116]) );
  LATCHX1 \decodedPacket_f_reg[1][115]  ( .CLK(n5876), .D(N9916), .Q(
        decodedPacket1_o[115]) );
  LATCHX1 \decodedPacket_f_reg[1][114]  ( .CLK(n5876), .D(N9915), .Q(
        decodedPacket1_o[114]) );
  LATCHX1 \decodedPacket_f_reg[1][113]  ( .CLK(n5876), .D(N9914), .Q(
        decodedPacket1_o[113]) );
  LATCHX1 \decodedPacket_f_reg[1][112]  ( .CLK(n5876), .D(N9913), .Q(
        decodedPacket1_o[112]) );
  LATCHX1 \decodedPacket_f_reg[1][111]  ( .CLK(n5876), .D(N9912), .Q(
        decodedPacket1_o[111]) );
  LATCHX1 \decodedPacket_f_reg[1][110]  ( .CLK(n5876), .D(N9911), .Q(
        decodedPacket1_o[110]) );
  LATCHX1 \decodedPacket_f_reg[1][109]  ( .CLK(n5876), .D(N9910), .Q(
        decodedPacket1_o[109]) );
  LATCHX1 \decodedPacket_f_reg[1][108]  ( .CLK(n5876), .D(N9909), .Q(
        decodedPacket1_o[108]) );
  LATCHX1 \decodedPacket_f_reg[1][107]  ( .CLK(n5875), .D(N9908), .Q(
        decodedPacket1_o[107]) );
  LATCHX1 \decodedPacket_f_reg[1][106]  ( .CLK(n5875), .D(N9907), .Q(
        decodedPacket1_o[106]) );
  LATCHX1 \decodedPacket_f_reg[1][105]  ( .CLK(n5875), .D(N9906), .Q(
        decodedPacket1_o[105]) );
  LATCHX1 \decodedPacket_f_reg[1][104]  ( .CLK(n5875), .D(N9905), .Q(
        decodedPacket1_o[104]) );
  LATCHX1 \decodedPacket_f_reg[1][103]  ( .CLK(n5875), .D(N9904), .Q(
        decodedPacket1_o[103]) );
  LATCHX1 \decodedPacket_f_reg[1][102]  ( .CLK(n5875), .D(N9903), .Q(
        decodedPacket1_o[102]) );
  LATCHX1 \decodedPacket_f_reg[1][101]  ( .CLK(n5875), .D(N9902), .Q(
        decodedPacket1_o[101]) );
  LATCHX1 \decodedPacket_f_reg[1][100]  ( .CLK(n5875), .D(N9901), .Q(
        decodedPacket1_o[100]) );
  LATCHX1 \decodedPacket_f_reg[1][99]  ( .CLK(n5875), .D(N9900), .Q(
        decodedPacket1_o[99]) );
  LATCHX1 \decodedPacket_f_reg[1][98]  ( .CLK(n5875), .D(N9898), .Q(
        decodedPacket1_o[98]) );
  LATCHX1 \decodedPacket_f_reg[1][97]  ( .CLK(n5875), .D(N9896), .Q(
        decodedPacket1_o[97]) );
  LATCHX1 \decodedPacket_f_reg[1][96]  ( .CLK(n5875), .D(N9895), .Q(
        decodedPacket1_o[96]) );
  LATCHX1 \decodedPacket_f_reg[1][95]  ( .CLK(n5874), .D(N9894), .Q(
        decodedPacket1_o[95]) );
  LATCHX1 \decodedPacket_f_reg[1][94]  ( .CLK(n5874), .D(N9893), .Q(
        decodedPacket1_o[94]) );
  LATCHX1 \decodedPacket_f_reg[1][93]  ( .CLK(n5874), .D(N9892), .Q(
        decodedPacket1_o[93]) );
  LATCHX1 \decodedPacket_f_reg[1][92]  ( .CLK(n5874), .D(N9891), .Q(
        decodedPacket1_o[92]) );
  LATCHX1 \decodedPacket_f_reg[1][91]  ( .CLK(n5874), .D(N9890), .Q(
        decodedPacket1_o[91]) );
  LATCHX1 \decodedPacket_f_reg[1][90]  ( .CLK(n5874), .D(N9889), .Q(
        decodedPacket1_o[90]) );
  LATCHX1 \decodedPacket_f_reg[1][89]  ( .CLK(n5874), .D(N9888), .Q(
        decodedPacket1_o[89]) );
  LATCHX1 \decodedPacket_f_reg[1][88]  ( .CLK(n5874), .D(N9887), .Q(
        decodedPacket1_o[88]) );
  LATCHX1 \decodedPacket_f_reg[1][87]  ( .CLK(n5874), .D(N9886), .Q(
        decodedPacket1_o[87]) );
  LATCHX1 \decodedPacket_f_reg[1][86]  ( .CLK(n5874), .D(N9885), .Q(
        decodedPacket1_o[86]) );
  LATCHX1 \decodedPacket_f_reg[1][85]  ( .CLK(n5874), .D(N9884), .Q(
        decodedPacket1_o[85]) );
  LATCHX1 \decodedPacket_f_reg[1][84]  ( .CLK(n5874), .D(N9883), .Q(
        decodedPacket1_o[84]) );
  LATCHX1 \decodedPacket_f_reg[1][83]  ( .CLK(n5873), .D(N9882), .Q(
        decodedPacket1_o[83]) );
  LATCHX1 \decodedPacket_f_reg[1][82]  ( .CLK(n5873), .D(N9881), .Q(
        decodedPacket1_o[82]) );
  LATCHX1 \decodedPacket_f_reg[1][81]  ( .CLK(n5873), .D(N9880), .Q(
        decodedPacket1_o[81]) );
  LATCHX1 \decodedPacket_f_reg[1][80]  ( .CLK(n5873), .D(N9879), .Q(
        decodedPacket1_o[80]) );
  LATCHX1 \decodedPacket_f_reg[1][79]  ( .CLK(n5873), .D(N9878), .Q(
        decodedPacket1_o[79]) );
  LATCHX1 \decodedPacket_f_reg[1][78]  ( .CLK(n5873), .D(N9877), .Q(
        decodedPacket1_o[78]) );
  LATCHX1 \decodedPacket_f_reg[1][77]  ( .CLK(n5873), .D(N9876), .Q(
        decodedPacket1_o[77]) );
  LATCHX1 \decodedPacket_f_reg[1][76]  ( .CLK(n5873), .D(N9875), .Q(
        decodedPacket1_o[76]) );
  LATCHX1 \decodedPacket_f_reg[1][75]  ( .CLK(n5873), .D(N9874), .Q(
        decodedPacket1_o[75]) );
  LATCHX1 \decodedPacket_f_reg[1][74]  ( .CLK(n5873), .D(N9873), .Q(
        decodedPacket1_o[74]) );
  LATCHX1 \decodedPacket_f_reg[1][73]  ( .CLK(n5873), .D(N9872), .Q(
        decodedPacket1_o[73]) );
  LATCHX1 \decodedPacket_f_reg[1][72]  ( .CLK(n5873), .D(N9871), .Q(
        decodedPacket1_o[72]) );
  LATCHX1 \decodedPacket_f_reg[1][71]  ( .CLK(n5872), .D(N9870), .Q(
        decodedPacket1_o[71]) );
  LATCHX1 \decodedPacket_f_reg[1][70]  ( .CLK(n5872), .D(N9869), .Q(
        decodedPacket1_o[70]) );
  LATCHX1 \decodedPacket_f_reg[1][69]  ( .CLK(n5872), .D(N9868), .Q(
        decodedPacket1_o[69]) );
  LATCHX1 \decodedPacket_f_reg[1][68]  ( .CLK(n5872), .D(N9867), .Q(
        decodedPacket1_o[68]) );
  LATCHX1 \decodedPacket_f_reg[1][67]  ( .CLK(n5872), .D(N9866), .Q(
        decodedPacket1_o[67]) );
  LATCHX1 \decodedPacket_f_reg[1][66]  ( .CLK(n5872), .D(N9865), .Q(
        decodedPacket1_o[66]) );
  LATCHX1 \decodedPacket_f_reg[1][65]  ( .CLK(n5872), .D(N9864), .Q(
        decodedPacket1_o[65]) );
  LATCHX1 \decodedPacket_f_reg[1][64]  ( .CLK(n5872), .D(N9863), .Q(
        decodedPacket1_o[64]) );
  LATCHX1 \decodedPacket_f_reg[1][63]  ( .CLK(n5872), .D(N9862), .Q(
        decodedPacket1_o[63]) );
  LATCHX1 \decodedPacket_f_reg[1][62]  ( .CLK(n5872), .D(N9861), .Q(
        decodedPacket1_o[62]) );
  LATCHX1 \decodedPacket_f_reg[1][61]  ( .CLK(n5872), .D(N9860), .Q(
        decodedPacket1_o[61]) );
  LATCHX1 \decodedPacket_f_reg[1][60]  ( .CLK(n5872), .D(N9859), .Q(
        decodedPacket1_o[60]) );
  LATCHX1 \decodedPacket_f_reg[1][59]  ( .CLK(n5871), .D(N9858), .Q(
        decodedPacket1_o[59]) );
  LATCHX1 \decodedPacket_f_reg[1][58]  ( .CLK(n5871), .D(N9857), .Q(
        decodedPacket1_o[58]) );
  LATCHX1 \decodedPacket_f_reg[1][57]  ( .CLK(n5871), .D(N9856), .Q(
        decodedPacket1_o[57]) );
  LATCHX1 \decodedPacket_f_reg[1][56]  ( .CLK(n5871), .D(N9855), .Q(
        decodedPacket1_o[56]) );
  LATCHX1 \decodedPacket_f_reg[1][55]  ( .CLK(n5871), .D(N9854), .Q(
        decodedPacket1_o[55]) );
  LATCHX1 \decodedPacket_f_reg[1][54]  ( .CLK(n5871), .D(N9853), .Q(
        decodedPacket1_o[54]) );
  LATCHX1 \decodedPacket_f_reg[1][53]  ( .CLK(n5871), .D(N9852), .Q(
        decodedPacket1_o[53]) );
  LATCHX1 \decodedPacket_f_reg[1][52]  ( .CLK(n5871), .D(N9851), .Q(
        decodedPacket1_o[52]) );
  LATCHX1 \decodedPacket_f_reg[1][51]  ( .CLK(n5871), .D(N9850), .Q(
        decodedPacket1_o[51]) );
  LATCHX1 \decodedPacket_f_reg[1][50]  ( .CLK(n5871), .D(N9849), .Q(
        decodedPacket1_o[50]) );
  LATCHX1 \decodedPacket_f_reg[1][49]  ( .CLK(n5871), .D(N9848), .Q(
        decodedPacket1_o[49]) );
  LATCHX1 \decodedPacket_f_reg[1][48]  ( .CLK(n5871), .D(N9846), .Q(
        decodedPacket1_o[48]) );
  LATCHX1 \decodedPacket_f_reg[1][47]  ( .CLK(n5870), .D(N9845), .Q(
        decodedPacket1_o[47]) );
  LATCHX1 \decodedPacket_f_reg[1][46]  ( .CLK(n5870), .D(N9844), .Q(
        decodedPacket1_o[46]) );
  LATCHX1 \decodedPacket_f_reg[1][45]  ( .CLK(n5870), .D(N9843), .Q(
        decodedPacket1_o[45]) );
  LATCHX1 \decodedPacket_f_reg[1][44]  ( .CLK(n5870), .D(N9842), .Q(
        decodedPacket1_o[44]) );
  LATCHX1 \decodedPacket_f_reg[1][43]  ( .CLK(n5870), .D(N9841), .Q(
        decodedPacket1_o[43]) );
  LATCHX1 \decodedPacket_f_reg[1][42]  ( .CLK(n5870), .D(N9840), .Q(
        decodedPacket1_o[42]) );
  LATCHX1 \decodedPacket_f_reg[1][41]  ( .CLK(n5870), .D(N9839), .Q(
        decodedPacket1_o[41]) );
  LATCHX1 \decodedPacket_f_reg[1][40]  ( .CLK(n5870), .D(N9838), .Q(
        decodedPacket1_o[40]) );
  LATCHX1 \decodedPacket_f_reg[1][39]  ( .CLK(n5870), .D(N9837), .Q(
        decodedPacket1_o[39]) );
  LATCHX1 \decodedPacket_f_reg[1][38]  ( .CLK(n5870), .D(N9836), .Q(
        decodedPacket1_o[38]) );
  LATCHX1 \decodedPacket_f_reg[1][37]  ( .CLK(n5870), .D(N9835), .Q(
        decodedPacket1_o[37]) );
  LATCHX1 \decodedPacket_f_reg[1][36]  ( .CLK(n5870), .D(N9834), .Q(
        decodedPacket1_o[36]) );
  LATCHX1 \decodedPacket_f_reg[1][35]  ( .CLK(n5869), .D(N9833), .Q(
        decodedPacket1_o[35]) );
  LATCHX1 \decodedPacket_f_reg[1][34]  ( .CLK(n5869), .D(N9832), .Q(
        decodedPacket1_o[34]) );
  LATCHX1 \decodedPacket_f_reg[1][33]  ( .CLK(n5869), .D(N9831), .Q(
        decodedPacket1_o[33]) );
  LATCHX1 \decodedPacket_f_reg[1][32]  ( .CLK(n5869), .D(N9830), .Q(
        decodedPacket1_o[32]) );
  LATCHX1 \decodedPacket_f_reg[1][31]  ( .CLK(n5869), .D(N9829), .Q(
        decodedPacket1_o[31]) );
  LATCHX1 \decodedPacket_f_reg[1][30]  ( .CLK(n5869), .D(N9828), .Q(
        decodedPacket1_o[30]) );
  LATCHX1 \decodedPacket_f_reg[1][29]  ( .CLK(n5869), .D(N9827), .Q(
        decodedPacket1_o[29]) );
  LATCHX1 \decodedPacket_f_reg[1][28]  ( .CLK(n5869), .D(N9826), .Q(
        decodedPacket1_o[28]) );
  LATCHX1 \decodedPacket_f_reg[1][27]  ( .CLK(n5869), .D(N9825), .Q(
        decodedPacket1_o[27]) );
  LATCHX1 \decodedPacket_f_reg[1][26]  ( .CLK(n5869), .D(N9824), .Q(
        decodedPacket1_o[26]) );
  LATCHX1 \decodedPacket_f_reg[1][25]  ( .CLK(n5869), .D(N9823), .Q(
        decodedPacket1_o[25]) );
  LATCHX1 \decodedPacket_f_reg[1][24]  ( .CLK(n5869), .D(N9822), .Q(
        decodedPacket1_o[24]) );
  LATCHX1 \decodedPacket_f_reg[1][23]  ( .CLK(n5868), .D(N9821), .Q(
        decodedPacket1_o[23]) );
  LATCHX1 \decodedPacket_f_reg[1][22]  ( .CLK(n5868), .D(N9820), .Q(
        decodedPacket1_o[22]) );
  LATCHX1 \decodedPacket_f_reg[1][21]  ( .CLK(n5868), .D(N9819), .Q(
        decodedPacket1_o[21]) );
  LATCHX1 \decodedPacket_f_reg[1][20]  ( .CLK(n5868), .D(N9818), .Q(
        decodedPacket1_o[20]) );
  LATCHX1 \decodedPacket_f_reg[1][19]  ( .CLK(n5868), .D(N9817), .Q(
        decodedPacket1_o[19]) );
  LATCHX1 \decodedPacket_f_reg[1][18]  ( .CLK(n5868), .D(N9816), .Q(
        decodedPacket1_o[18]) );
  LATCHX1 \decodedPacket_f_reg[1][17]  ( .CLK(n5868), .D(N9815), .Q(
        decodedPacket1_o[17]) );
  LATCHX1 \decodedPacket_f_reg[1][16]  ( .CLK(n5868), .D(N9814), .Q(
        decodedPacket1_o[16]) );
  LATCHX1 \decodedPacket_f_reg[1][15]  ( .CLK(n5868), .D(N9813), .Q(
        decodedPacket1_o[15]) );
  LATCHX1 \decodedPacket_f_reg[1][14]  ( .CLK(n5868), .D(N9812), .Q(
        decodedPacket1_o[14]) );
  LATCHX1 \decodedPacket_f_reg[1][13]  ( .CLK(n5868), .D(N9811), .Q(
        decodedPacket1_o[13]) );
  LATCHX1 \decodedPacket_f_reg[1][12]  ( .CLK(n5868), .D(N9810), .Q(
        decodedPacket1_o[12]) );
  LATCHX1 \decodedPacket_f_reg[1][11]  ( .CLK(n5867), .D(N9809), .Q(
        decodedPacket1_o[11]) );
  LATCHX1 \decodedPacket_f_reg[1][10]  ( .CLK(n5867), .D(N9808), .Q(
        decodedPacket1_o[10]) );
  LATCHX1 \decodedPacket_f_reg[1][9]  ( .CLK(n5867), .D(N9807), .Q(
        decodedPacket1_o[9]) );
  LATCHX1 \decodedPacket_f_reg[1][8]  ( .CLK(n5867), .D(N9806), .Q(
        decodedPacket1_o[8]) );
  LATCHX1 \decodedPacket_f_reg[1][7]  ( .CLK(n5867), .D(N9805), .Q(
        decodedPacket1_o[7]) );
  LATCHX1 \decodedPacket_f_reg[1][6]  ( .CLK(n5867), .D(N9804), .Q(
        decodedPacket1_o[6]) );
  LATCHX1 \decodedPacket_f_reg[1][5]  ( .CLK(n5867), .D(N9803), .Q(
        decodedPacket1_o[5]) );
  LATCHX1 \decodedPacket_f_reg[1][4]  ( .CLK(n5867), .D(N9802), .Q(
        decodedPacket1_o[4]) );
  LATCHX1 \decodedPacket_f_reg[1][3]  ( .CLK(n5867), .D(N9801), .Q(
        decodedPacket1_o[3]) );
  LATCHX1 \decodedPacket_f_reg[1][2]  ( .CLK(n5867), .D(N9800), .Q(
        decodedPacket1_o[2]) );
  LATCHX1 \decodedPacket_f_reg[1][1]  ( .CLK(n5867), .D(N9799), .Q(
        decodedPacket1_o[1]) );
  LATCHX1 \decodedPacket_f_reg[1][0]  ( .CLK(n5867), .D(N9798), .Q(
        decodedPacket1_o[0]) );
  LATCHX1 \decodedPacket_f_reg[0][121]  ( .CLK(n5861), .D(N9792), .Q(
        decodedPacket0_o[121]) );
  LATCHX1 \decodedPacket_f_reg[0][120]  ( .CLK(n5862), .D(N9791), .Q(
        decodedPacket0_o[120]) );
  LATCHX1 \decodedPacket_f_reg[0][119]  ( .CLK(n5866), .D(N9790), .Q(
        decodedPacket0_o[119]) );
  LATCHX1 \decodedPacket_f_reg[0][118]  ( .CLK(n5866), .D(N9789), .Q(
        decodedPacket0_o[118]) );
  LATCHX1 \decodedPacket_f_reg[0][117]  ( .CLK(n5866), .D(N9788), .Q(
        decodedPacket0_o[117]) );
  LATCHX1 \decodedPacket_f_reg[0][116]  ( .CLK(n5866), .D(N9787), .Q(
        decodedPacket0_o[116]) );
  LATCHX1 \decodedPacket_f_reg[0][115]  ( .CLK(n5866), .D(N9786), .Q(
        decodedPacket0_o[115]) );
  LATCHX1 \decodedPacket_f_reg[0][114]  ( .CLK(n5866), .D(N9785), .Q(
        decodedPacket0_o[114]) );
  LATCHX1 \decodedPacket_f_reg[0][113]  ( .CLK(n5866), .D(N9784), .Q(
        decodedPacket0_o[113]) );
  LATCHX1 \decodedPacket_f_reg[0][112]  ( .CLK(n5866), .D(N9783), .Q(
        decodedPacket0_o[112]) );
  LATCHX1 \decodedPacket_f_reg[0][111]  ( .CLK(n5866), .D(N9782), .Q(
        decodedPacket0_o[111]) );
  LATCHX1 \decodedPacket_f_reg[0][110]  ( .CLK(n5866), .D(N9781), .Q(
        decodedPacket0_o[110]) );
  LATCHX1 \decodedPacket_f_reg[0][109]  ( .CLK(n5866), .D(N9780), .Q(
        decodedPacket0_o[109]) );
  LATCHX1 \decodedPacket_f_reg[0][108]  ( .CLK(n5866), .D(N9779), .Q(
        decodedPacket0_o[108]) );
  LATCHX1 \decodedPacket_f_reg[0][107]  ( .CLK(n5865), .D(N9778), .Q(
        decodedPacket0_o[107]) );
  LATCHX1 \decodedPacket_f_reg[0][106]  ( .CLK(n5865), .D(N9777), .Q(
        decodedPacket0_o[106]) );
  LATCHX1 \decodedPacket_f_reg[0][105]  ( .CLK(n5865), .D(N9776), .Q(
        decodedPacket0_o[105]) );
  LATCHX1 \decodedPacket_f_reg[0][104]  ( .CLK(n5865), .D(N9775), .Q(
        decodedPacket0_o[104]) );
  LATCHX1 \decodedPacket_f_reg[0][103]  ( .CLK(n5865), .D(N9774), .Q(
        decodedPacket0_o[103]) );
  LATCHX1 \decodedPacket_f_reg[0][102]  ( .CLK(n5865), .D(N9773), .Q(
        decodedPacket0_o[102]) );
  LATCHX1 \decodedPacket_f_reg[0][101]  ( .CLK(n5865), .D(N9772), .Q(
        decodedPacket0_o[101]) );
  LATCHX1 \decodedPacket_f_reg[0][100]  ( .CLK(n5865), .D(N9771), .Q(
        decodedPacket0_o[100]) );
  LATCHX1 \decodedPacket_f_reg[0][99]  ( .CLK(n5865), .D(N9770), .Q(
        decodedPacket0_o[99]) );
  LATCHX1 \decodedPacket_f_reg[0][98]  ( .CLK(n5865), .D(N9769), .Q(
        decodedPacket0_o[98]) );
  LATCHX1 \decodedPacket_f_reg[0][97]  ( .CLK(n5865), .D(N9768), .Q(
        decodedPacket0_o[97]) );
  LATCHX1 \decodedPacket_f_reg[0][96]  ( .CLK(n5865), .D(N9766), .Q(
        decodedPacket0_o[96]) );
  LATCHX1 \decodedPacket_f_reg[0][95]  ( .CLK(n5864), .D(N9765), .Q(
        decodedPacket0_o[95]) );
  LATCHX1 \decodedPacket_f_reg[0][94]  ( .CLK(n5864), .D(N9764), .Q(
        decodedPacket0_o[94]) );
  LATCHX1 \decodedPacket_f_reg[0][93]  ( .CLK(n5864), .D(N9763), .Q(
        decodedPacket0_o[93]) );
  LATCHX1 \decodedPacket_f_reg[0][92]  ( .CLK(n5864), .D(N9762), .Q(
        decodedPacket0_o[92]) );
  LATCHX1 \decodedPacket_f_reg[0][91]  ( .CLK(n5864), .D(N9761), .Q(
        decodedPacket0_o[91]) );
  LATCHX1 \decodedPacket_f_reg[0][90]  ( .CLK(n5864), .D(N9760), .Q(
        decodedPacket0_o[90]) );
  LATCHX1 \decodedPacket_f_reg[0][89]  ( .CLK(n5864), .D(N9759), .Q(
        decodedPacket0_o[89]) );
  LATCHX1 \decodedPacket_f_reg[0][88]  ( .CLK(n5864), .D(N9758), .Q(
        decodedPacket0_o[88]) );
  LATCHX1 \decodedPacket_f_reg[0][87]  ( .CLK(n5864), .D(N9757), .Q(
        decodedPacket0_o[87]) );
  LATCHX1 \decodedPacket_f_reg[0][86]  ( .CLK(n5864), .D(N9756), .Q(
        decodedPacket0_o[86]) );
  LATCHX1 \decodedPacket_f_reg[0][85]  ( .CLK(n5864), .D(N9755), .Q(
        decodedPacket0_o[85]) );
  LATCHX1 \decodedPacket_f_reg[0][84]  ( .CLK(n5864), .D(N9754), .Q(
        decodedPacket0_o[84]) );
  LATCHX1 \decodedPacket_f_reg[0][83]  ( .CLK(n5863), .D(N9753), .Q(
        decodedPacket0_o[83]) );
  LATCHX1 \decodedPacket_f_reg[0][82]  ( .CLK(n5863), .D(N9752), .Q(
        decodedPacket0_o[82]) );
  LATCHX1 \decodedPacket_f_reg[0][81]  ( .CLK(n5863), .D(N9751), .Q(
        decodedPacket0_o[81]) );
  LATCHX1 \decodedPacket_f_reg[0][80]  ( .CLK(n5863), .D(N9750), .Q(
        decodedPacket0_o[80]) );
  LATCHX1 \decodedPacket_f_reg[0][79]  ( .CLK(n5863), .D(N9749), .Q(
        decodedPacket0_o[79]) );
  LATCHX1 \decodedPacket_f_reg[0][78]  ( .CLK(n5863), .D(N9748), .Q(
        decodedPacket0_o[78]) );
  LATCHX1 \decodedPacket_f_reg[0][77]  ( .CLK(n5863), .D(N9747), .Q(
        decodedPacket0_o[77]) );
  LATCHX1 \decodedPacket_f_reg[0][76]  ( .CLK(n5863), .D(N9746), .Q(
        decodedPacket0_o[76]) );
  LATCHX1 \decodedPacket_f_reg[0][75]  ( .CLK(n5863), .D(N9745), .Q(
        decodedPacket0_o[75]) );
  LATCHX1 \decodedPacket_f_reg[0][74]  ( .CLK(n5863), .D(N9744), .Q(
        decodedPacket0_o[74]) );
  LATCHX1 \decodedPacket_f_reg[0][73]  ( .CLK(n5863), .D(N9743), .Q(
        decodedPacket0_o[73]) );
  LATCHX1 \decodedPacket_f_reg[0][72]  ( .CLK(n5863), .D(N9742), .Q(
        decodedPacket0_o[72]) );
  LATCHX1 \decodedPacket_f_reg[0][71]  ( .CLK(n5862), .D(N9741), .Q(
        decodedPacket0_o[71]) );
  LATCHX1 \decodedPacket_f_reg[0][70]  ( .CLK(n5862), .D(N9740), .Q(
        decodedPacket0_o[70]) );
  LATCHX1 \decodedPacket_f_reg[0][69]  ( .CLK(n5862), .D(N9739), .Q(
        decodedPacket0_o[69]) );
  LATCHX1 \decodedPacket_f_reg[0][68]  ( .CLK(n5862), .D(N9738), .Q(
        decodedPacket0_o[68]) );
  LATCHX1 \decodedPacket_f_reg[0][67]  ( .CLK(n5862), .D(N9737), .Q(
        decodedPacket0_o[67]) );
  LATCHX1 \decodedPacket_f_reg[0][66]  ( .CLK(n5862), .D(N9736), .Q(
        decodedPacket0_o[66]) );
  LATCHX1 \decodedPacket_f_reg[0][65]  ( .CLK(n5862), .D(N9735), .Q(
        decodedPacket0_o[65]) );
  LATCHX1 \decodedPacket_f_reg[0][64]  ( .CLK(n5862), .D(N9734), .Q(
        decodedPacket0_o[64]) );
  LATCHX1 \decodedPacket_f_reg[0][63]  ( .CLK(n5862), .D(N9733), .Q(
        decodedPacket0_o[63]) );
  LATCHX1 \decodedPacket_f_reg[0][62]  ( .CLK(n5862), .D(N9732), .Q(
        decodedPacket0_o[62]) );
  LATCHX1 \decodedPacket_f_reg[0][61]  ( .CLK(n5862), .D(N9731), .Q(
        decodedPacket0_o[61]) );
  LATCHX1 \decodedPacket_f_reg[0][60]  ( .CLK(n5862), .D(N9730), .Q(
        decodedPacket0_o[60]) );
  LATCHX1 \decodedPacket_f_reg[0][59]  ( .CLK(n5861), .D(N9729), .Q(
        decodedPacket0_o[59]) );
  LATCHX1 \decodedPacket_f_reg[0][58]  ( .CLK(n5861), .D(N9728), .Q(
        decodedPacket0_o[58]) );
  LATCHX1 \decodedPacket_f_reg[0][57]  ( .CLK(n5861), .D(N9727), .Q(
        decodedPacket0_o[57]) );
  LATCHX1 \decodedPacket_f_reg[0][56]  ( .CLK(n5861), .D(N9726), .Q(
        decodedPacket0_o[56]) );
  LATCHX1 \decodedPacket_f_reg[0][55]  ( .CLK(n5861), .D(N9725), .Q(
        decodedPacket0_o[55]) );
  LATCHX1 \decodedPacket_f_reg[0][54]  ( .CLK(n5861), .D(N9724), .Q(
        decodedPacket0_o[54]) );
  LATCHX1 \decodedPacket_f_reg[0][53]  ( .CLK(n5861), .D(N9723), .Q(
        decodedPacket0_o[53]) );
  LATCHX1 \decodedPacket_f_reg[0][52]  ( .CLK(n5861), .D(N9722), .Q(
        decodedPacket0_o[52]) );
  LATCHX1 \decodedPacket_f_reg[0][51]  ( .CLK(n5861), .D(N9721), .Q(
        decodedPacket0_o[51]) );
  LATCHX1 \decodedPacket_f_reg[0][50]  ( .CLK(n5861), .D(N9720), .Q(
        decodedPacket0_o[50]) );
  LATCHX1 \decodedPacket_f_reg[0][49]  ( .CLK(n5861), .D(N9719), .Q(
        decodedPacket0_o[49]) );
  LATCHX1 \decodedPacket_f_reg[0][48]  ( .CLK(n5861), .D(N9718), .Q(
        decodedPacket0_o[48]) );
  LATCHX1 \decodedPacket_f_reg[0][47]  ( .CLK(n5860), .D(N9716), .Q(
        decodedPacket0_o[47]) );
  LATCHX1 \decodedPacket_f_reg[0][46]  ( .CLK(n5860), .D(N9715), .Q(
        decodedPacket0_o[46]) );
  LATCHX1 \decodedPacket_f_reg[0][45]  ( .CLK(n5860), .D(N9714), .Q(
        decodedPacket0_o[45]) );
  LATCHX1 \decodedPacket_f_reg[0][44]  ( .CLK(n5860), .D(N9713), .Q(
        decodedPacket0_o[44]) );
  LATCHX1 \decodedPacket_f_reg[0][43]  ( .CLK(n5860), .D(N9712), .Q(
        decodedPacket0_o[43]) );
  LATCHX1 \decodedPacket_f_reg[0][42]  ( .CLK(n5860), .D(N9711), .Q(
        decodedPacket0_o[42]) );
  LATCHX1 \decodedPacket_f_reg[0][41]  ( .CLK(n5860), .D(N9710), .Q(
        decodedPacket0_o[41]) );
  LATCHX1 \decodedPacket_f_reg[0][40]  ( .CLK(n5860), .D(N9709), .Q(
        decodedPacket0_o[40]) );
  LATCHX1 \decodedPacket_f_reg[0][39]  ( .CLK(n5860), .D(N9708), .Q(
        decodedPacket0_o[39]) );
  LATCHX1 \decodedPacket_f_reg[0][38]  ( .CLK(n5860), .D(N9707), .Q(
        decodedPacket0_o[38]) );
  LATCHX1 \decodedPacket_f_reg[0][37]  ( .CLK(n5860), .D(N9706), .Q(
        decodedPacket0_o[37]) );
  LATCHX1 \decodedPacket_f_reg[0][36]  ( .CLK(n5860), .D(N9705), .Q(
        decodedPacket0_o[36]) );
  LATCHX1 \decodedPacket_f_reg[0][35]  ( .CLK(n5859), .D(N9704), .Q(
        decodedPacket0_o[35]) );
  LATCHX1 \decodedPacket_f_reg[0][34]  ( .CLK(n5859), .D(N9703), .Q(
        decodedPacket0_o[34]) );
  LATCHX1 \decodedPacket_f_reg[0][33]  ( .CLK(n5859), .D(N9702), .Q(
        decodedPacket0_o[33]) );
  LATCHX1 \decodedPacket_f_reg[0][32]  ( .CLK(n5859), .D(N9701), .Q(
        decodedPacket0_o[32]) );
  LATCHX1 \decodedPacket_f_reg[0][31]  ( .CLK(n5859), .D(N9700), .Q(
        decodedPacket0_o[31]) );
  LATCHX1 \decodedPacket_f_reg[0][30]  ( .CLK(n5859), .D(N9699), .Q(
        decodedPacket0_o[30]) );
  LATCHX1 \decodedPacket_f_reg[0][29]  ( .CLK(n5859), .D(N9698), .Q(
        decodedPacket0_o[29]) );
  LATCHX1 \decodedPacket_f_reg[0][28]  ( .CLK(n5859), .D(N9697), .Q(
        decodedPacket0_o[28]) );
  LATCHX1 \decodedPacket_f_reg[0][27]  ( .CLK(n5859), .D(N9696), .Q(
        decodedPacket0_o[27]) );
  LATCHX1 \decodedPacket_f_reg[0][26]  ( .CLK(n5859), .D(N9695), .Q(
        decodedPacket0_o[26]) );
  LATCHX1 \decodedPacket_f_reg[0][25]  ( .CLK(n5859), .D(N9694), .Q(
        decodedPacket0_o[25]) );
  LATCHX1 \decodedPacket_f_reg[0][24]  ( .CLK(n5859), .D(N9693), .Q(
        decodedPacket0_o[24]) );
  LATCHX1 \decodedPacket_f_reg[0][23]  ( .CLK(n5858), .D(N9692), .Q(
        decodedPacket0_o[23]) );
  LATCHX1 \decodedPacket_f_reg[0][22]  ( .CLK(n5858), .D(N9691), .Q(
        decodedPacket0_o[22]) );
  LATCHX1 \decodedPacket_f_reg[0][21]  ( .CLK(n5858), .D(N9690), .Q(
        decodedPacket0_o[21]) );
  LATCHX1 \decodedPacket_f_reg[0][20]  ( .CLK(n5858), .D(N9689), .Q(
        decodedPacket0_o[20]) );
  LATCHX1 \decodedPacket_f_reg[0][19]  ( .CLK(n5858), .D(N9688), .Q(
        decodedPacket0_o[19]) );
  LATCHX1 \decodedPacket_f_reg[0][18]  ( .CLK(n5858), .D(N9687), .Q(
        decodedPacket0_o[18]) );
  LATCHX1 \decodedPacket_f_reg[0][17]  ( .CLK(n5858), .D(N9686), .Q(
        decodedPacket0_o[17]) );
  LATCHX1 \decodedPacket_f_reg[0][16]  ( .CLK(n5858), .D(N9685), .Q(
        decodedPacket0_o[16]) );
  LATCHX1 \decodedPacket_f_reg[0][15]  ( .CLK(n5858), .D(N9684), .Q(
        decodedPacket0_o[15]) );
  LATCHX1 \decodedPacket_f_reg[0][14]  ( .CLK(n5858), .D(N9683), .Q(
        decodedPacket0_o[14]) );
  LATCHX1 \decodedPacket_f_reg[0][13]  ( .CLK(n5858), .D(N9682), .Q(
        decodedPacket0_o[13]) );
  LATCHX1 \decodedPacket_f_reg[0][12]  ( .CLK(n5858), .D(N9681), .Q(
        decodedPacket0_o[12]) );
  LATCHX1 \decodedPacket_f_reg[0][11]  ( .CLK(n5857), .D(N9680), .Q(
        decodedPacket0_o[11]) );
  LATCHX1 \decodedPacket_f_reg[0][10]  ( .CLK(n5857), .D(N9679), .Q(
        decodedPacket0_o[10]) );
  LATCHX1 \decodedPacket_f_reg[0][9]  ( .CLK(n5857), .D(N9678), .Q(
        decodedPacket0_o[9]) );
  LATCHX1 \decodedPacket_f_reg[0][8]  ( .CLK(n5857), .D(N9677), .Q(
        decodedPacket0_o[8]) );
  LATCHX1 \decodedPacket_f_reg[0][7]  ( .CLK(n5857), .D(N9676), .Q(
        decodedPacket0_o[7]) );
  LATCHX1 \decodedPacket_f_reg[0][6]  ( .CLK(n5857), .D(N9675), .Q(
        decodedPacket0_o[6]) );
  LATCHX1 \decodedPacket_f_reg[0][5]  ( .CLK(n5857), .D(N9674), .Q(
        decodedPacket0_o[5]) );
  LATCHX1 \decodedPacket_f_reg[0][4]  ( .CLK(n5857), .D(N9673), .Q(
        decodedPacket0_o[4]) );
  LATCHX1 \decodedPacket_f_reg[0][3]  ( .CLK(n5857), .D(N9672), .Q(
        decodedPacket0_o[3]) );
  LATCHX1 \decodedPacket_f_reg[0][2]  ( .CLK(n5857), .D(N9671), .Q(
        decodedPacket0_o[2]) );
  LATCHX1 \decodedPacket_f_reg[0][1]  ( .CLK(n5857), .D(N9670), .Q(
        decodedPacket0_o[1]) );
  LATCHX1 \decodedPacket_f_reg[0][0]  ( .CLK(n5857), .D(N9669), .Q(
        decodedPacket0_o[0]) );
  OAI22X1 U868 ( .IN1(n5845), .IN2(n825), .IN3(n5849), .IN4(n6350), .QN(N9999)
         );
  OA22X1 U869 ( .IN1(n5826), .IN2(n827), .IN3(n5825), .IN4(n6351), .Q(n825) );
  OA22X1 U870 ( .IN1(n5812), .IN2(n6196), .IN3(n5818), .IN4(n830), .Q(n827) );
  OA22X1 U871 ( .IN1(n5790), .IN2(n831), .IN3(n5806), .IN4(n6197), .Q(n830) );
  OA22X1 U872 ( .IN1(n5777), .IN2(n6042), .IN3(n5779), .IN4(n6043), .Q(n831)
         );
  OAI22X1 U873 ( .IN1(n5845), .IN2(n834), .IN3(n5852), .IN4(n6395), .QN(N9998)
         );
  OA22X1 U874 ( .IN1(n5826), .IN2(n835), .IN3(n5838), .IN4(n6392), .Q(n834) );
  OA22X1 U875 ( .IN1(n5810), .IN2(n6243), .IN3(n5816), .IN4(n836), .Q(n835) );
  OA22X1 U876 ( .IN1(n5790), .IN2(n837), .IN3(n5800), .IN4(n6238), .Q(n836) );
  OA22X1 U877 ( .IN1(n5775), .IN2(n6089), .IN3(n5781), .IN4(n6084), .Q(n837)
         );
  OAI22X1 U878 ( .IN1(n5845), .IN2(n838), .IN3(n5848), .IN4(n6423), .QN(N9997)
         );
  OA22X1 U879 ( .IN1(n5826), .IN2(n839), .IN3(n5825), .IN4(n6423), .Q(n838) );
  OA22X1 U880 ( .IN1(n5810), .IN2(n6269), .IN3(n5819), .IN4(n840), .Q(n839) );
  OA22X1 U881 ( .IN1(n5790), .IN2(n841), .IN3(n5807), .IN4(n6269), .Q(n840) );
  OA22X1 U882 ( .IN1(n5775), .IN2(n6115), .IN3(n5781), .IN4(n6115), .Q(n841)
         );
  OAI22X1 U883 ( .IN1(n5845), .IN2(n842), .IN3(n5853), .IN4(n6424), .QN(N9996)
         );
  OA22X1 U884 ( .IN1(n5826), .IN2(n843), .IN3(n5841), .IN4(n6424), .Q(n842) );
  OA22X1 U885 ( .IN1(n5810), .IN2(n6270), .IN3(n5816), .IN4(n844), .Q(n843) );
  OA22X1 U886 ( .IN1(n5790), .IN2(n845), .IN3(n5801), .IN4(n6270), .Q(n844) );
  OA22X1 U887 ( .IN1(n5775), .IN2(n6116), .IN3(n5782), .IN4(n6116), .Q(n845)
         );
  OAI22X1 U888 ( .IN1(n5845), .IN2(n846), .IN3(n5848), .IN4(n6425), .QN(N9995)
         );
  OA22X1 U889 ( .IN1(n5826), .IN2(n847), .IN3(n5840), .IN4(n6425), .Q(n846) );
  OA22X1 U890 ( .IN1(n5810), .IN2(n6271), .IN3(n5814), .IN4(n848), .Q(n847) );
  OA22X1 U891 ( .IN1(n5790), .IN2(n849), .IN3(n5805), .IN4(n6271), .Q(n848) );
  OA22X1 U892 ( .IN1(n5775), .IN2(n6117), .IN3(n5779), .IN4(n6117), .Q(n849)
         );
  OAI22X1 U893 ( .IN1(n5845), .IN2(n850), .IN3(n5848), .IN4(n6426), .QN(N9994)
         );
  OA22X1 U894 ( .IN1(n5826), .IN2(n851), .IN3(n5842), .IN4(n6426), .Q(n850) );
  OA22X1 U895 ( .IN1(n5811), .IN2(n6272), .IN3(n5814), .IN4(n852), .Q(n851) );
  OA22X1 U896 ( .IN1(n5790), .IN2(n853), .IN3(n5787), .IN4(n6272), .Q(n852) );
  OA22X1 U897 ( .IN1(n5775), .IN2(n6118), .IN3(n5779), .IN4(n6118), .Q(n853)
         );
  OAI22X1 U898 ( .IN1(n5845), .IN2(n854), .IN3(n5848), .IN4(n6427), .QN(N9993)
         );
  OA22X1 U899 ( .IN1(n5826), .IN2(n855), .IN3(n5842), .IN4(n6427), .Q(n854) );
  OA22X1 U900 ( .IN1(n5811), .IN2(n6273), .IN3(n5814), .IN4(n856), .Q(n855) );
  OA22X1 U901 ( .IN1(n5790), .IN2(n857), .IN3(n5788), .IN4(n6273), .Q(n856) );
  OA22X1 U902 ( .IN1(n5776), .IN2(n6119), .IN3(n5779), .IN4(n6119), .Q(n857)
         );
  OAI22X1 U903 ( .IN1(n5846), .IN2(n858), .IN3(n5848), .IN4(n6428), .QN(N9992)
         );
  OA22X1 U904 ( .IN1(n5826), .IN2(n859), .IN3(n5825), .IN4(n6428), .Q(n858) );
  OA22X1 U905 ( .IN1(n5811), .IN2(n6274), .IN3(n5814), .IN4(n860), .Q(n859) );
  OA22X1 U906 ( .IN1(n5790), .IN2(n861), .IN3(n5789), .IN4(n6274), .Q(n860) );
  OA22X1 U907 ( .IN1(n5776), .IN2(n6120), .IN3(n5779), .IN4(n6120), .Q(n861)
         );
  OAI22X1 U908 ( .IN1(n5846), .IN2(n862), .IN3(n5848), .IN4(n6429), .QN(N9991)
         );
  OA22X1 U909 ( .IN1(n5826), .IN2(n863), .IN3(n5825), .IN4(n6429), .Q(n862) );
  OA22X1 U910 ( .IN1(n5811), .IN2(n6275), .IN3(n5814), .IN4(n864), .Q(n863) );
  OA22X1 U911 ( .IN1(n5790), .IN2(n865), .IN3(n5802), .IN4(n6275), .Q(n864) );
  OA22X1 U912 ( .IN1(n5776), .IN2(n6121), .IN3(n5779), .IN4(n6121), .Q(n865)
         );
  OAI22X1 U913 ( .IN1(n5846), .IN2(n866), .IN3(n5849), .IN4(n6430), .QN(N9990)
         );
  OA22X1 U914 ( .IN1(n5826), .IN2(n867), .IN3(n5837), .IN4(n6430), .Q(n866) );
  OA22X1 U915 ( .IN1(n5811), .IN2(n6276), .IN3(n5815), .IN4(n868), .Q(n867) );
  OA22X1 U916 ( .IN1(n5790), .IN2(n869), .IN3(n5803), .IN4(n6276), .Q(n868) );
  OA22X1 U917 ( .IN1(n5776), .IN2(n6122), .IN3(n5780), .IN4(n6122), .Q(n869)
         );
  OAI22X1 U918 ( .IN1(n5846), .IN2(n870), .IN3(n5849), .IN4(n6431), .QN(N9989)
         );
  OA22X1 U919 ( .IN1(n5826), .IN2(n871), .IN3(n5839), .IN4(n6431), .Q(n870) );
  OA22X1 U920 ( .IN1(n5811), .IN2(n6277), .IN3(n5819), .IN4(n872), .Q(n871) );
  OA22X1 U921 ( .IN1(n5790), .IN2(n873), .IN3(n5803), .IN4(n6277), .Q(n872) );
  OA22X1 U922 ( .IN1(n5776), .IN2(n6123), .IN3(n5780), .IN4(n6123), .Q(n873)
         );
  OAI22X1 U923 ( .IN1(n5846), .IN2(n874), .IN3(n5849), .IN4(n6432), .QN(N9988)
         );
  OA22X1 U924 ( .IN1(n5826), .IN2(n875), .IN3(n5823), .IN4(n6432), .Q(n874) );
  OA22X1 U925 ( .IN1(n5811), .IN2(n6278), .IN3(n5819), .IN4(n876), .Q(n875) );
  OA22X1 U926 ( .IN1(n5790), .IN2(n877), .IN3(n5804), .IN4(n6278), .Q(n876) );
  OA22X1 U927 ( .IN1(n5776), .IN2(n6124), .IN3(n5780), .IN4(n6124), .Q(n877)
         );
  OAI22X1 U928 ( .IN1(n5846), .IN2(n878), .IN3(n5849), .IN4(n6433), .QN(N9987)
         );
  OA22X1 U929 ( .IN1(n5827), .IN2(n879), .IN3(n5824), .IN4(n6433), .Q(n878) );
  OA22X1 U930 ( .IN1(n5811), .IN2(n6279), .IN3(n5819), .IN4(n880), .Q(n879) );
  OA22X1 U931 ( .IN1(n5791), .IN2(n881), .IN3(n5803), .IN4(n6279), .Q(n880) );
  OA22X1 U932 ( .IN1(n5776), .IN2(n6125), .IN3(n5780), .IN4(n6125), .Q(n881)
         );
  OAI22X1 U933 ( .IN1(n5846), .IN2(n882), .IN3(n5849), .IN4(n6434), .QN(N9986)
         );
  OA22X1 U934 ( .IN1(n5827), .IN2(n883), .IN3(n5825), .IN4(n6434), .Q(n882) );
  OA22X1 U935 ( .IN1(n5811), .IN2(n6280), .IN3(n5816), .IN4(n884), .Q(n883) );
  OA22X1 U936 ( .IN1(n5791), .IN2(n885), .IN3(n5806), .IN4(n6280), .Q(n884) );
  OA22X1 U937 ( .IN1(n5776), .IN2(n6126), .IN3(n5780), .IN4(n6126), .Q(n885)
         );
  OAI22X1 U938 ( .IN1(n5846), .IN2(n886), .IN3(n5850), .IN4(n6435), .QN(N9985)
         );
  OA22X1 U939 ( .IN1(n5827), .IN2(n887), .IN3(n5824), .IN4(n6435), .Q(n886) );
  OA22X1 U940 ( .IN1(n5811), .IN2(n6281), .IN3(n5817), .IN4(n888), .Q(n887) );
  OA22X1 U941 ( .IN1(n5791), .IN2(n889), .IN3(n5788), .IN4(n6281), .Q(n888) );
  OA22X1 U942 ( .IN1(n5776), .IN2(n6127), .IN3(n5784), .IN4(n6127), .Q(n889)
         );
  OAI22X1 U943 ( .IN1(n5846), .IN2(n890), .IN3(n5850), .IN4(n6436), .QN(N9984)
         );
  OA22X1 U944 ( .IN1(n5827), .IN2(n891), .IN3(n5836), .IN4(n6436), .Q(n890) );
  OA22X1 U945 ( .IN1(n5811), .IN2(n6282), .IN3(n5819), .IN4(n892), .Q(n891) );
  OA22X1 U946 ( .IN1(n5791), .IN2(n893), .IN3(n5789), .IN4(n6282), .Q(n892) );
  OA22X1 U947 ( .IN1(n5776), .IN2(n6128), .IN3(n5786), .IN4(n6128), .Q(n893)
         );
  OAI22X1 U948 ( .IN1(n5846), .IN2(n894), .IN3(n5850), .IN4(n6437), .QN(N9983)
         );
  OA22X1 U949 ( .IN1(n5827), .IN2(n895), .IN3(n5825), .IN4(n6437), .Q(n894) );
  OA22X1 U950 ( .IN1(n5811), .IN2(n6283), .IN3(n5816), .IN4(n896), .Q(n895) );
  OA22X1 U951 ( .IN1(n5791), .IN2(n897), .IN3(n5800), .IN4(n6283), .Q(n896) );
  OA22X1 U952 ( .IN1(n5776), .IN2(n6129), .IN3(n5783), .IN4(n6129), .Q(n897)
         );
  OAI22X1 U953 ( .IN1(n5846), .IN2(n898), .IN3(n5850), .IN4(n6438), .QN(N9982)
         );
  OA22X1 U954 ( .IN1(n5827), .IN2(n899), .IN3(n5837), .IN4(n6438), .Q(n898) );
  OA22X1 U955 ( .IN1(n5811), .IN2(n6284), .IN3(n5817), .IN4(n900), .Q(n899) );
  OA22X1 U956 ( .IN1(n5791), .IN2(n901), .IN3(n5787), .IN4(n6284), .Q(n900) );
  OA22X1 U957 ( .IN1(n5776), .IN2(n6130), .IN3(n5783), .IN4(n6130), .Q(n901)
         );
  OAI22X1 U958 ( .IN1(n5846), .IN2(n902), .IN3(n5850), .IN4(n6439), .QN(N9981)
         );
  OA22X1 U959 ( .IN1(n5827), .IN2(n903), .IN3(n5839), .IN4(n6439), .Q(n902) );
  OA22X1 U960 ( .IN1(n5811), .IN2(n6285), .IN3(n5820), .IN4(n904), .Q(n903) );
  OA22X1 U961 ( .IN1(n5791), .IN2(n905), .IN3(n5807), .IN4(n6285), .Q(n904) );
  OA22X1 U962 ( .IN1(n5776), .IN2(n6131), .IN3(n5783), .IN4(n6131), .Q(n905)
         );
  OAI22X1 U963 ( .IN1(n5846), .IN2(n906), .IN3(n826), .IN4(n6440), .QN(N9980)
         );
  OA22X1 U964 ( .IN1(n5827), .IN2(n907), .IN3(n5840), .IN4(n6440), .Q(n906) );
  OA22X1 U965 ( .IN1(n5811), .IN2(n6286), .IN3(n5817), .IN4(n908), .Q(n907) );
  OA22X1 U966 ( .IN1(n5791), .IN2(n909), .IN3(n5787), .IN4(n6286), .Q(n908) );
  OA22X1 U967 ( .IN1(n5776), .IN2(n6132), .IN3(n5785), .IN4(n6132), .Q(n909)
         );
  OAI22X1 U968 ( .IN1(n5846), .IN2(n910), .IN3(n826), .IN4(n6441), .QN(N9979)
         );
  OA22X1 U969 ( .IN1(n5827), .IN2(n911), .IN3(n5838), .IN4(n6441), .Q(n910) );
  OA22X1 U970 ( .IN1(n5811), .IN2(n6287), .IN3(n5820), .IN4(n912), .Q(n911) );
  OA22X1 U971 ( .IN1(n5791), .IN2(n913), .IN3(n5789), .IN4(n6287), .Q(n912) );
  OA22X1 U972 ( .IN1(n5776), .IN2(n6133), .IN3(n5784), .IN4(n6133), .Q(n913)
         );
  OAI22X1 U973 ( .IN1(n5846), .IN2(n914), .IN3(n826), .IN4(n6442), .QN(N9978)
         );
  OA22X1 U974 ( .IN1(n5827), .IN2(n915), .IN3(n5824), .IN4(n6442), .Q(n914) );
  OA22X1 U975 ( .IN1(n5811), .IN2(n6288), .IN3(n5814), .IN4(n916), .Q(n915) );
  OA22X1 U976 ( .IN1(n5791), .IN2(n917), .IN3(n5788), .IN4(n6288), .Q(n916) );
  OA22X1 U977 ( .IN1(n5776), .IN2(n6134), .IN3(n5786), .IN4(n6134), .Q(n917)
         );
  OAI22X1 U978 ( .IN1(n5846), .IN2(n918), .IN3(n826), .IN4(n6443), .QN(N9976)
         );
  OA22X1 U979 ( .IN1(n5827), .IN2(n919), .IN3(n5841), .IN4(n6443), .Q(n918) );
  OA22X1 U980 ( .IN1(n5811), .IN2(n6289), .IN3(n5815), .IN4(n920), .Q(n919) );
  OA22X1 U981 ( .IN1(n5791), .IN2(n921), .IN3(n5802), .IN4(n6289), .Q(n920) );
  OA22X1 U982 ( .IN1(n5776), .IN2(n6135), .IN3(n5782), .IN4(n6135), .Q(n921)
         );
  OAI22X1 U983 ( .IN1(n5846), .IN2(n922), .IN3(n826), .IN4(n6444), .QN(N9975)
         );
  OA22X1 U984 ( .IN1(n5827), .IN2(n923), .IN3(n5840), .IN4(n6444), .Q(n922) );
  OA22X1 U985 ( .IN1(n5811), .IN2(n6290), .IN3(n5818), .IN4(n924), .Q(n923) );
  OA22X1 U986 ( .IN1(n5791), .IN2(n925), .IN3(n5807), .IN4(n6290), .Q(n924) );
  OA22X1 U987 ( .IN1(n5776), .IN2(n6136), .IN3(n5783), .IN4(n6136), .Q(n925)
         );
  OAI22X1 U988 ( .IN1(n5846), .IN2(n926), .IN3(n5853), .IN4(n6445), .QN(N9974)
         );
  OA22X1 U989 ( .IN1(n5828), .IN2(n927), .IN3(n5837), .IN4(n6445), .Q(n926) );
  OA22X1 U990 ( .IN1(n5811), .IN2(n6291), .IN3(n5815), .IN4(n928), .Q(n927) );
  OA22X1 U991 ( .IN1(n5792), .IN2(n929), .IN3(n5805), .IN4(n6291), .Q(n928) );
  OA22X1 U992 ( .IN1(n5776), .IN2(n6137), .IN3(n5781), .IN4(n6137), .Q(n929)
         );
  OAI22X1 U993 ( .IN1(n5846), .IN2(n930), .IN3(n5850), .IN4(n6446), .QN(N9973)
         );
  OA22X1 U994 ( .IN1(n5828), .IN2(n931), .IN3(n5836), .IN4(n6446), .Q(n930) );
  OA22X1 U995 ( .IN1(n5811), .IN2(n6292), .IN3(n5815), .IN4(n932), .Q(n931) );
  OA22X1 U996 ( .IN1(n5792), .IN2(n933), .IN3(n5802), .IN4(n6292), .Q(n932) );
  OA22X1 U997 ( .IN1(n5776), .IN2(n6138), .IN3(n5781), .IN4(n6138), .Q(n933)
         );
  OAI22X1 U998 ( .IN1(n5846), .IN2(n934), .IN3(n5848), .IN4(n6447), .QN(N9972)
         );
  OA22X1 U999 ( .IN1(n5828), .IN2(n935), .IN3(n5836), .IN4(n6447), .Q(n934) );
  OA22X1 U1000 ( .IN1(n5811), .IN2(n6293), .IN3(n5815), .IN4(n936), .Q(n935)
         );
  OA22X1 U1001 ( .IN1(n5792), .IN2(n937), .IN3(n5803), .IN4(n6293), .Q(n936)
         );
  OA22X1 U1002 ( .IN1(n5776), .IN2(n6139), .IN3(n5781), .IN4(n6139), .Q(n937)
         );
  OAI22X1 U1003 ( .IN1(n5846), .IN2(n938), .IN3(n5852), .IN4(n6448), .QN(N9971) );
  OA22X1 U1004 ( .IN1(n5828), .IN2(n939), .IN3(n5824), .IN4(n6448), .Q(n938)
         );
  OA22X1 U1005 ( .IN1(n5811), .IN2(n6294), .IN3(n5815), .IN4(n940), .Q(n939)
         );
  OA22X1 U1006 ( .IN1(n5792), .IN2(n941), .IN3(n5804), .IN4(n6294), .Q(n940)
         );
  OA22X1 U1007 ( .IN1(n5776), .IN2(n6140), .IN3(n5781), .IN4(n6140), .Q(n941)
         );
  OAI22X1 U1008 ( .IN1(n5846), .IN2(n942), .IN3(n826), .IN4(n6449), .QN(N9970)
         );
  OA22X1 U1009 ( .IN1(n5828), .IN2(n943), .IN3(n5842), .IN4(n6449), .Q(n942)
         );
  OA22X1 U1010 ( .IN1(n5811), .IN2(n6295), .IN3(n5815), .IN4(n944), .Q(n943)
         );
  OA22X1 U1011 ( .IN1(n5792), .IN2(n945), .IN3(n5800), .IN4(n6295), .Q(n944)
         );
  OA22X1 U1012 ( .IN1(n5776), .IN2(n6141), .IN3(n5781), .IN4(n6141), .Q(n945)
         );
  OAI22X1 U1013 ( .IN1(n5846), .IN2(n946), .IN3(n5852), .IN4(n6450), .QN(N9969) );
  OA22X1 U1014 ( .IN1(n5828), .IN2(n947), .IN3(n5822), .IN4(n6450), .Q(n946)
         );
  OA22X1 U1015 ( .IN1(n5811), .IN2(n6296), .IN3(n5820), .IN4(n948), .Q(n947)
         );
  OA22X1 U1016 ( .IN1(n5792), .IN2(n949), .IN3(n5800), .IN4(n6296), .Q(n948)
         );
  OA22X1 U1017 ( .IN1(n5776), .IN2(n6142), .IN3(n5781), .IN4(n6142), .Q(n949)
         );
  OAI22X1 U1018 ( .IN1(n5846), .IN2(n950), .IN3(n5849), .IN4(n6451), .QN(N9968) );
  OA22X1 U1019 ( .IN1(n5828), .IN2(n951), .IN3(n5823), .IN4(n6451), .Q(n950)
         );
  OA22X1 U1020 ( .IN1(n5811), .IN2(n6297), .IN3(n5814), .IN4(n952), .Q(n951)
         );
  OA22X1 U1021 ( .IN1(n5792), .IN2(n953), .IN3(n5787), .IN4(n6297), .Q(n952)
         );
  OA22X1 U1022 ( .IN1(n5776), .IN2(n6143), .IN3(n5779), .IN4(n6143), .Q(n953)
         );
  OAI22X1 U1023 ( .IN1(n5846), .IN2(n954), .IN3(n826), .IN4(n6452), .QN(N9967)
         );
  OA22X1 U1024 ( .IN1(n5828), .IN2(n955), .IN3(n5839), .IN4(n6452), .Q(n954)
         );
  OA22X1 U1025 ( .IN1(n5811), .IN2(n6298), .IN3(n5815), .IN4(n956), .Q(n955)
         );
  OA22X1 U1026 ( .IN1(n5792), .IN2(n957), .IN3(n5789), .IN4(n6298), .Q(n956)
         );
  OA22X1 U1027 ( .IN1(n5776), .IN2(n6144), .IN3(n5785), .IN4(n6144), .Q(n957)
         );
  OAI22X1 U1028 ( .IN1(n5846), .IN2(n958), .IN3(n5850), .IN4(n6453), .QN(N9966) );
  OA22X1 U1029 ( .IN1(n5828), .IN2(n959), .IN3(n5838), .IN4(n6453), .Q(n958)
         );
  OA22X1 U1030 ( .IN1(n5811), .IN2(n6299), .IN3(n5818), .IN4(n960), .Q(n959)
         );
  OA22X1 U1031 ( .IN1(n5792), .IN2(n961), .IN3(n5788), .IN4(n6299), .Q(n960)
         );
  OA22X1 U1032 ( .IN1(n5776), .IN2(n6145), .IN3(n5784), .IN4(n6145), .Q(n961)
         );
  OAI22X1 U1033 ( .IN1(n5846), .IN2(n962), .IN3(n5852), .IN4(n6454), .QN(N9965) );
  OA22X1 U1034 ( .IN1(n5828), .IN2(n963), .IN3(n5839), .IN4(n6454), .Q(n962)
         );
  OA22X1 U1035 ( .IN1(n5811), .IN2(n6300), .IN3(n5821), .IN4(n964), .Q(n963)
         );
  OA22X1 U1036 ( .IN1(n5792), .IN2(n965), .IN3(n5801), .IN4(n6300), .Q(n964)
         );
  OA22X1 U1037 ( .IN1(n5776), .IN2(n6146), .IN3(n5786), .IN4(n6146), .Q(n965)
         );
  OA22X1 U1039 ( .IN1(n5828), .IN2(n967), .IN3(n5841), .IN4(n6320), .Q(n966)
         );
  OA22X1 U1044 ( .IN1(n5828), .IN2(n971), .IN3(n5825), .IN4(n6321), .Q(n970)
         );
  OA22X1 U1049 ( .IN1(n5829), .IN2(n975), .IN3(n5823), .IN4(n6322), .Q(n974)
         );
  OA22X1 U1054 ( .IN1(n5829), .IN2(n979), .IN3(n5840), .IN4(n6323), .Q(n978)
         );
  OA22X1 U1059 ( .IN1(n5829), .IN2(n983), .IN3(n5841), .IN4(n6324), .Q(n982)
         );
  OA22X1 U1064 ( .IN1(n5829), .IN2(n987), .IN3(n5842), .IN4(n6325), .Q(n986)
         );
  OA22X1 U1069 ( .IN1(n5829), .IN2(n991), .IN3(n5836), .IN4(n6326), .Q(n990)
         );
  OA22X1 U1074 ( .IN1(n5829), .IN2(n995), .IN3(n5823), .IN4(n6327), .Q(n994)
         );
  OA22X1 U1079 ( .IN1(n5829), .IN2(n999), .IN3(n5824), .IN4(n6328), .Q(n998)
         );
  OA22X1 U1084 ( .IN1(n5829), .IN2(n1003), .IN3(n5842), .IN4(n6329), .Q(n1002)
         );
  OA22X1 U1089 ( .IN1(n5829), .IN2(n1007), .IN3(n5839), .IN4(n6330), .Q(n1006)
         );
  OA22X1 U1094 ( .IN1(n5829), .IN2(n1011), .IN3(n5837), .IN4(n6331), .Q(n1010)
         );
  OA22X1 U1099 ( .IN1(n5829), .IN2(n1015), .IN3(n5838), .IN4(n6332), .Q(n1014)
         );
  OA22X1 U1104 ( .IN1(n5829), .IN2(n1019), .IN3(n5836), .IN4(n6333), .Q(n1018)
         );
  OA22X1 U1109 ( .IN1(n5830), .IN2(n1023), .IN3(n5836), .IN4(n6334), .Q(n1022)
         );
  OA22X1 U1114 ( .IN1(n5830), .IN2(n1027), .IN3(n5836), .IN4(n6335), .Q(n1026)
         );
  OA22X1 U1119 ( .IN1(n5830), .IN2(n1031), .IN3(n5836), .IN4(n6336), .Q(n1030)
         );
  OA22X1 U1124 ( .IN1(n5830), .IN2(n1035), .IN3(n5836), .IN4(n6337), .Q(n1034)
         );
  OA22X1 U1129 ( .IN1(n5830), .IN2(n1039), .IN3(n5841), .IN4(n6338), .Q(n1038)
         );
  OA22X1 U1134 ( .IN1(n5830), .IN2(n1043), .IN3(n5824), .IN4(n6339), .Q(n1042)
         );
  OA22X1 U1139 ( .IN1(n5830), .IN2(n1047), .IN3(n5839), .IN4(n6340), .Q(n1046)
         );
  OA22X1 U1144 ( .IN1(n5830), .IN2(n1051), .IN3(n5825), .IN4(n6341), .Q(n1050)
         );
  OA22X1 U1149 ( .IN1(n5830), .IN2(n1055), .IN3(n5822), .IN4(n6342), .Q(n1054)
         );
  OA22X1 U1154 ( .IN1(n5830), .IN2(n1059), .IN3(n5839), .IN4(n6343), .Q(n1058)
         );
  OA22X1 U1159 ( .IN1(n5830), .IN2(n1063), .IN3(n5822), .IN4(n6344), .Q(n1062)
         );
  OA22X1 U1164 ( .IN1(n5830), .IN2(n1067), .IN3(n5823), .IN4(n6345), .Q(n1066)
         );
  OA22X1 U1169 ( .IN1(n5831), .IN2(n1071), .IN3(n5824), .IN4(n6346), .Q(n1070)
         );
  OA22X1 U1174 ( .IN1(n5831), .IN2(n1075), .IN3(n5837), .IN4(n6315), .Q(n1074)
         );
  OA22X1 U1179 ( .IN1(n5831), .IN2(n1079), .IN3(n5837), .IN4(n6316), .Q(n1078)
         );
  OA22X1 U1184 ( .IN1(n5831), .IN2(n1083), .IN3(n5837), .IN4(n6317), .Q(n1082)
         );
  OA22X1 U1189 ( .IN1(n5831), .IN2(n1087), .IN3(n5837), .IN4(n6318), .Q(n1086)
         );
  OA22X1 U1194 ( .IN1(n5831), .IN2(n1091), .IN3(n5837), .IN4(n6319), .Q(n1090)
         );
  OAI22X1 U1198 ( .IN1(n5846), .IN2(n1094), .IN3(n5851), .IN4(n6455), .QN(
        N9932) );
  OA22X1 U1199 ( .IN1(n5831), .IN2(n1095), .IN3(n5838), .IN4(n6455), .Q(n1094)
         );
  OA22X1 U1200 ( .IN1(n5811), .IN2(n6301), .IN3(n5816), .IN4(n1096), .Q(n1095)
         );
  OA22X1 U1201 ( .IN1(n5795), .IN2(n1097), .IN3(n5800), .IN4(n6301), .Q(n1096)
         );
  OA22X1 U1202 ( .IN1(n5776), .IN2(n6147), .IN3(n5782), .IN4(n6147), .Q(n1097)
         );
  OAI22X1 U1203 ( .IN1(n5846), .IN2(n1098), .IN3(n5851), .IN4(n6456), .QN(
        N9931) );
  OA22X1 U1204 ( .IN1(n5831), .IN2(n1099), .IN3(n5838), .IN4(n6456), .Q(n1098)
         );
  OA22X1 U1205 ( .IN1(n5811), .IN2(n6302), .IN3(n5816), .IN4(n1100), .Q(n1099)
         );
  OA22X1 U1206 ( .IN1(n5795), .IN2(n1101), .IN3(n5800), .IN4(n6302), .Q(n1100)
         );
  OA22X1 U1207 ( .IN1(n5776), .IN2(n6148), .IN3(n5782), .IN4(n6148), .Q(n1101)
         );
  OAI22X1 U1208 ( .IN1(n5846), .IN2(n1102), .IN3(n5851), .IN4(n6457), .QN(
        N9930) );
  OA22X1 U1209 ( .IN1(n5831), .IN2(n1103), .IN3(n5838), .IN4(n6457), .Q(n1102)
         );
  OA22X1 U1210 ( .IN1(n5812), .IN2(n6303), .IN3(n5816), .IN4(n1104), .Q(n1103)
         );
  OA22X1 U1211 ( .IN1(n5795), .IN2(n1105), .IN3(n5801), .IN4(n6303), .Q(n1104)
         );
  OA22X1 U1212 ( .IN1(n5776), .IN2(n6149), .IN3(n5782), .IN4(n6149), .Q(n1105)
         );
  OAI22X1 U1213 ( .IN1(n5846), .IN2(n1106), .IN3(n5851), .IN4(n6458), .QN(
        N9929) );
  OA22X1 U1214 ( .IN1(n5831), .IN2(n1107), .IN3(n5838), .IN4(n6458), .Q(n1106)
         );
  OA22X1 U1215 ( .IN1(n5812), .IN2(n6304), .IN3(n5816), .IN4(n1108), .Q(n1107)
         );
  OA22X1 U1216 ( .IN1(n5795), .IN2(n1109), .IN3(n5801), .IN4(n6304), .Q(n1108)
         );
  OA22X1 U1217 ( .IN1(n5777), .IN2(n6150), .IN3(n5782), .IN4(n6150), .Q(n1109)
         );
  OAI22X1 U1218 ( .IN1(n5846), .IN2(n1110), .IN3(n5851), .IN4(n6459), .QN(
        N9928) );
  OA22X1 U1219 ( .IN1(n5831), .IN2(n1111), .IN3(n5838), .IN4(n6459), .Q(n1110)
         );
  OA22X1 U1220 ( .IN1(n5812), .IN2(n6305), .IN3(n5816), .IN4(n1112), .Q(n1111)
         );
  OA22X1 U1221 ( .IN1(n5795), .IN2(n1113), .IN3(n5801), .IN4(n6305), .Q(n1112)
         );
  OA22X1 U1222 ( .IN1(n5777), .IN2(n6151), .IN3(n5782), .IN4(n6151), .Q(n1113)
         );
  OA22X1 U1248 ( .IN1(n5743), .IN2(n5856), .IN3(n5753), .IN4(n1141), .Q(n1140)
         );
  OAI22X1 U1253 ( .IN1(n5770), .IN2(n6384), .IN3(n5763), .IN4(n1145), .QN(
        N9921) );
  OA22X1 U1254 ( .IN1(n5741), .IN2(n6349), .IN3(n5756), .IN4(n1146), .Q(n1145)
         );
  OA22X1 U1255 ( .IN1(n5740), .IN2(n1147), .IN3(n5731), .IN4(n6230), .Q(n1146)
         );
  OA22X1 U1256 ( .IN1(n5708), .IN2(n6195), .IN3(n5717), .IN4(n1148), .Q(n1147)
         );
  OA22X1 U1257 ( .IN1(n5707), .IN2(n1149), .IN3(n5700), .IN4(n6076), .Q(n1148)
         );
  AOI22X1 U1258 ( .IN1(n5695), .IN2(\decodedPacket[2][120] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][120] ), .QN(n1149) );
  OAI22X1 U1259 ( .IN1(n5766), .IN2(n6376), .IN3(n5763), .IN4(n1150), .QN(
        N9920) );
  OA22X1 U1260 ( .IN1(n5741), .IN2(n6348), .IN3(n5757), .IN4(n1151), .Q(n1150)
         );
  OA22X1 U1261 ( .IN1(n5740), .IN2(n1152), .IN3(n5729), .IN4(n6222), .Q(n1151)
         );
  OA22X1 U1262 ( .IN1(n5708), .IN2(n6194), .IN3(n5718), .IN4(n1153), .Q(n1152)
         );
  OA22X1 U1263 ( .IN1(n5707), .IN2(n1154), .IN3(n5698), .IN4(n6068), .Q(n1153)
         );
  AOI22X1 U1264 ( .IN1(n5695), .IN2(\decodedPacket[2][119] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][119] ), .QN(n1154) );
  OAI22X1 U1265 ( .IN1(n5766), .IN2(n6372), .IN3(n5763), .IN4(n1155), .QN(
        N9919) );
  OA22X1 U1266 ( .IN1(n5741), .IN2(n6374), .IN3(n5750), .IN4(n1156), .Q(n1155)
         );
  OA22X1 U1267 ( .IN1(n5740), .IN2(n1157), .IN3(n5729), .IN4(n6219), .Q(n1156)
         );
  OA22X1 U1268 ( .IN1(n5708), .IN2(n6220), .IN3(n5721), .IN4(n1158), .Q(n1157)
         );
  OA22X1 U1269 ( .IN1(n5707), .IN2(n1159), .IN3(n5698), .IN4(n6064), .Q(n1158)
         );
  AOI22X1 U1270 ( .IN1(n5695), .IN2(\decodedPacket[2][118] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][118] ), .QN(n1159) );
  OA22X1 U1272 ( .IN1(n5741), .IN2(n6371), .IN3(n5753), .IN4(n1161), .Q(n1160)
         );
  OAI22X1 U1277 ( .IN1(n5766), .IN2(n6373), .IN3(n5763), .IN4(n1165), .QN(
        N9917) );
  OA22X1 U1278 ( .IN1(n5741), .IN2(n6370), .IN3(n5759), .IN4(n1166), .Q(n1165)
         );
  OA22X1 U1279 ( .IN1(n5740), .IN2(n1167), .IN3(n5729), .IN4(n6219), .Q(n1166)
         );
  OA22X1 U1280 ( .IN1(n5708), .IN2(n6216), .IN3(n5725), .IN4(n1168), .Q(n1167)
         );
  OA22X1 U1281 ( .IN1(n5707), .IN2(n1169), .IN3(n5698), .IN4(n6065), .Q(n1168)
         );
  AOI22X1 U1282 ( .IN1(n5695), .IN2(\decodedPacket[2][116] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][116] ), .QN(n1169) );
  OAI22X1 U1283 ( .IN1(n5766), .IN2(n6396), .IN3(n5763), .IN4(n1170), .QN(
        N9916) );
  OA22X1 U1284 ( .IN1(n5741), .IN2(n6347), .IN3(n5755), .IN4(n1171), .Q(n1170)
         );
  OA22X1 U1285 ( .IN1(n5739), .IN2(n1172), .IN3(n5729), .IN4(n6245), .Q(n1171)
         );
  OA22X1 U1286 ( .IN1(n5708), .IN2(n6193), .IN3(n5717), .IN4(n1173), .Q(n1172)
         );
  OA22X1 U1287 ( .IN1(n5707), .IN2(n1174), .IN3(n5698), .IN4(n6091), .Q(n1173)
         );
  AOI22X1 U1288 ( .IN1(n5695), .IN2(\decodedPacket[2][115] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][115] ), .QN(n1174) );
  OAI22X1 U1289 ( .IN1(n5766), .IN2(n5967), .IN3(n5763), .IN4(n1175), .QN(
        N9915) );
  OA22X1 U1290 ( .IN1(n5741), .IN2(n6369), .IN3(n5750), .IN4(n1176), .Q(n1175)
         );
  OA22X1 U1291 ( .IN1(n5739), .IN2(n1177), .IN3(n5729), .IN4(n5952), .Q(n1176)
         );
  OA22X1 U1292 ( .IN1(n5708), .IN2(n6215), .IN3(n5717), .IN4(n1178), .Q(n1177)
         );
  OA22X1 U1293 ( .IN1(n5707), .IN2(n1179), .IN3(n5698), .IN4(n5937), .Q(n1178)
         );
  AOI22X1 U1294 ( .IN1(n5695), .IN2(\decodedPacket[2][114] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][114] ), .QN(n1179) );
  OAI22X1 U1295 ( .IN1(n5766), .IN2(n5968), .IN3(n5764), .IN4(n1180), .QN(
        N9914) );
  OA22X1 U1296 ( .IN1(n5741), .IN2(n6368), .IN3(n5751), .IN4(n1181), .Q(n1180)
         );
  OA22X1 U1297 ( .IN1(n5739), .IN2(n1182), .IN3(n5730), .IN4(n5953), .Q(n1181)
         );
  OA22X1 U1298 ( .IN1(n5708), .IN2(n6214), .IN3(n5717), .IN4(n1183), .Q(n1182)
         );
  OA22X1 U1299 ( .IN1(n5707), .IN2(n1184), .IN3(n5698), .IN4(n5938), .Q(n1183)
         );
  AOI22X1 U1300 ( .IN1(n5695), .IN2(\decodedPacket[2][113] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][113] ), .QN(n1184) );
  OAI22X1 U1301 ( .IN1(n5766), .IN2(n5969), .IN3(n5764), .IN4(n1185), .QN(
        N9913) );
  OA22X1 U1302 ( .IN1(n5741), .IN2(n6367), .IN3(n5752), .IN4(n1186), .Q(n1185)
         );
  OA22X1 U1303 ( .IN1(n5739), .IN2(n1187), .IN3(n5730), .IN4(n5954), .Q(n1186)
         );
  OA22X1 U1304 ( .IN1(n5708), .IN2(n6213), .IN3(n5717), .IN4(n1188), .Q(n1187)
         );
  OA22X1 U1305 ( .IN1(n5707), .IN2(n1189), .IN3(n5699), .IN4(n5939), .Q(n1188)
         );
  AOI22X1 U1306 ( .IN1(n5695), .IN2(\decodedPacket[2][112] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][112] ), .QN(n1189) );
  OAI22X1 U1307 ( .IN1(n5767), .IN2(n5970), .IN3(n5764), .IN4(n1190), .QN(
        N9912) );
  OA22X1 U1308 ( .IN1(n5741), .IN2(n6366), .IN3(n5760), .IN4(n1191), .Q(n1190)
         );
  OA22X1 U1309 ( .IN1(n5739), .IN2(n1192), .IN3(n5730), .IN4(n5955), .Q(n1191)
         );
  OA22X1 U1310 ( .IN1(n5708), .IN2(n6212), .IN3(n5717), .IN4(n1193), .Q(n1192)
         );
  OA22X1 U1311 ( .IN1(n5707), .IN2(n1194), .IN3(n5699), .IN4(n5940), .Q(n1193)
         );
  AOI22X1 U1312 ( .IN1(n5695), .IN2(\decodedPacket[2][111] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][111] ), .QN(n1194) );
  OAI22X1 U1313 ( .IN1(n5767), .IN2(n5971), .IN3(n5764), .IN4(n1195), .QN(
        N9911) );
  OA22X1 U1314 ( .IN1(n5741), .IN2(n6365), .IN3(n5758), .IN4(n1196), .Q(n1195)
         );
  OA22X1 U1315 ( .IN1(n5739), .IN2(n1197), .IN3(n5730), .IN4(n5956), .Q(n1196)
         );
  OA22X1 U1316 ( .IN1(n5708), .IN2(n6211), .IN3(n5718), .IN4(n1198), .Q(n1197)
         );
  OA22X1 U1317 ( .IN1(n5707), .IN2(n1199), .IN3(n5699), .IN4(n5941), .Q(n1198)
         );
  AOI22X1 U1318 ( .IN1(n5695), .IN2(\decodedPacket[2][110] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][110] ), .QN(n1199) );
  OAI22X1 U1319 ( .IN1(n5767), .IN2(n5972), .IN3(n5764), .IN4(n1200), .QN(
        N9910) );
  OA22X1 U1320 ( .IN1(n5741), .IN2(n6364), .IN3(n5759), .IN4(n1201), .Q(n1200)
         );
  OA22X1 U1321 ( .IN1(n5739), .IN2(n1202), .IN3(n5730), .IN4(n5957), .Q(n1201)
         );
  OA22X1 U1322 ( .IN1(n5708), .IN2(n6210), .IN3(n5718), .IN4(n1203), .Q(n1202)
         );
  OA22X1 U1323 ( .IN1(n5707), .IN2(n1204), .IN3(n5699), .IN4(n5942), .Q(n1203)
         );
  AOI22X1 U1324 ( .IN1(n5695), .IN2(\decodedPacket[2][109] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][109] ), .QN(n1204) );
  OAI22X1 U1325 ( .IN1(n5767), .IN2(n5973), .IN3(n5764), .IN4(n1205), .QN(
        N9909) );
  OA22X1 U1326 ( .IN1(n5742), .IN2(n6363), .IN3(n5760), .IN4(n1206), .Q(n1205)
         );
  OA22X1 U1327 ( .IN1(n5739), .IN2(n1207), .IN3(n5730), .IN4(n5958), .Q(n1206)
         );
  OA22X1 U1328 ( .IN1(n5709), .IN2(n6209), .IN3(n5718), .IN4(n1208), .Q(n1207)
         );
  OA22X1 U1329 ( .IN1(n5706), .IN2(n1209), .IN3(n5699), .IN4(n5943), .Q(n1208)
         );
  AOI22X1 U1330 ( .IN1(n5695), .IN2(\decodedPacket[2][108] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][108] ), .QN(n1209) );
  OAI22X1 U1331 ( .IN1(n5767), .IN2(n5974), .IN3(n5764), .IN4(n1210), .QN(
        N9908) );
  OA22X1 U1332 ( .IN1(n5742), .IN2(n6362), .IN3(n5756), .IN4(n1211), .Q(n1210)
         );
  OA22X1 U1333 ( .IN1(n5739), .IN2(n1212), .IN3(n5730), .IN4(n5959), .Q(n1211)
         );
  OA22X1 U1334 ( .IN1(n5709), .IN2(n6208), .IN3(n5718), .IN4(n1213), .Q(n1212)
         );
  OA22X1 U1335 ( .IN1(n5705), .IN2(n1214), .IN3(n5699), .IN4(n5944), .Q(n1213)
         );
  AOI22X1 U1336 ( .IN1(n5695), .IN2(\decodedPacket[2][107] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][107] ), .QN(n1214) );
  OAI22X1 U1337 ( .IN1(n5767), .IN2(n5975), .IN3(n5764), .IN4(n1215), .QN(
        N9907) );
  OA22X1 U1338 ( .IN1(n5742), .IN2(n6308), .IN3(n5757), .IN4(n1216), .Q(n1215)
         );
  OA22X1 U1339 ( .IN1(n5739), .IN2(n1217), .IN3(n5730), .IN4(n5960), .Q(n1216)
         );
  OA22X1 U1340 ( .IN1(n5709), .IN2(n6154), .IN3(n5718), .IN4(n1218), .Q(n1217)
         );
  OA22X1 U1341 ( .IN1(n5704), .IN2(n1219), .IN3(n5699), .IN4(n5945), .Q(n1218)
         );
  AOI22X1 U1342 ( .IN1(n5695), .IN2(\decodedPacket[2][106] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][106] ), .QN(n1219) );
  OAI22X1 U1343 ( .IN1(n5767), .IN2(n5976), .IN3(n5764), .IN4(n1220), .QN(
        N9906) );
  OA22X1 U1344 ( .IN1(n5742), .IN2(n6309), .IN3(n5758), .IN4(n1221), .Q(n1220)
         );
  OA22X1 U1345 ( .IN1(n5739), .IN2(n1222), .IN3(n5730), .IN4(n5961), .Q(n1221)
         );
  OA22X1 U1346 ( .IN1(n5709), .IN2(n6155), .IN3(n5718), .IN4(n1223), .Q(n1222)
         );
  OA22X1 U1347 ( .IN1(n5706), .IN2(n1224), .IN3(n5699), .IN4(n5946), .Q(n1223)
         );
  AOI22X1 U1348 ( .IN1(n5695), .IN2(\decodedPacket[2][105] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][105] ), .QN(n1224) );
  OAI22X1 U1349 ( .IN1(n5767), .IN2(n5977), .IN3(n5764), .IN4(n1225), .QN(
        N9905) );
  OA22X1 U1350 ( .IN1(n5742), .IN2(n6310), .IN3(n5759), .IN4(n1226), .Q(n1225)
         );
  OA22X1 U1351 ( .IN1(n5739), .IN2(n1227), .IN3(n5730), .IN4(n5962), .Q(n1226)
         );
  OA22X1 U1352 ( .IN1(n5709), .IN2(n6156), .IN3(n5720), .IN4(n1228), .Q(n1227)
         );
  OA22X1 U1353 ( .IN1(n5706), .IN2(n1229), .IN3(n5699), .IN4(n5947), .Q(n1228)
         );
  AOI22X1 U1354 ( .IN1(n5695), .IN2(\decodedPacket[2][104] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][104] ), .QN(n1229) );
  OAI22X1 U1355 ( .IN1(n5767), .IN2(n5978), .IN3(n5764), .IN4(n1230), .QN(
        N9904) );
  OA22X1 U1356 ( .IN1(n5742), .IN2(n6311), .IN3(n5760), .IN4(n1231), .Q(n1230)
         );
  OA22X1 U1357 ( .IN1(n5738), .IN2(n1232), .IN3(n5730), .IN4(n5963), .Q(n1231)
         );
  OA22X1 U1358 ( .IN1(n5709), .IN2(n6157), .IN3(n5721), .IN4(n1233), .Q(n1232)
         );
  OA22X1 U1359 ( .IN1(n5706), .IN2(n1234), .IN3(n5699), .IN4(n5948), .Q(n1233)
         );
  AOI22X1 U1360 ( .IN1(n5695), .IN2(\decodedPacket[2][103] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][103] ), .QN(n1234) );
  OAI22X1 U1361 ( .IN1(n5767), .IN2(n5979), .IN3(n5764), .IN4(n1235), .QN(
        N9903) );
  OA22X1 U1362 ( .IN1(n5742), .IN2(n6312), .IN3(n5753), .IN4(n1236), .Q(n1235)
         );
  OA22X1 U1363 ( .IN1(n5738), .IN2(n1237), .IN3(n5730), .IN4(n5964), .Q(n1236)
         );
  OA22X1 U1364 ( .IN1(n5709), .IN2(n6158), .IN3(n5724), .IN4(n1238), .Q(n1237)
         );
  OA22X1 U1365 ( .IN1(n5706), .IN2(n1239), .IN3(n5699), .IN4(n5949), .Q(n1238)
         );
  AOI22X1 U1366 ( .IN1(n5695), .IN2(\decodedPacket[2][102] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][102] ), .QN(n1239) );
  OAI22X1 U1367 ( .IN1(n5767), .IN2(n5980), .IN3(n5764), .IN4(n1240), .QN(
        N9902) );
  OA22X1 U1368 ( .IN1(n5742), .IN2(n6313), .IN3(n5750), .IN4(n1241), .Q(n1240)
         );
  OA22X1 U1369 ( .IN1(n5738), .IN2(n1242), .IN3(n5730), .IN4(n5965), .Q(n1241)
         );
  OA22X1 U1370 ( .IN1(n5709), .IN2(n6159), .IN3(n5722), .IN4(n1243), .Q(n1242)
         );
  OA22X1 U1371 ( .IN1(n5706), .IN2(n1244), .IN3(n5699), .IN4(n5950), .Q(n1243)
         );
  AOI22X1 U1372 ( .IN1(n5695), .IN2(\decodedPacket[2][101] ), .IN3(n5683), 
        .IN4(\decodedPacket[1][101] ), .QN(n1244) );
  OAI22X1 U1373 ( .IN1(n5767), .IN2(n5981), .IN3(n5764), .IN4(n1245), .QN(
        N9901) );
  OA22X1 U1374 ( .IN1(n5742), .IN2(n6314), .IN3(n5759), .IN4(n1246), .Q(n1245)
         );
  OA22X1 U1375 ( .IN1(n5738), .IN2(n1247), .IN3(n5730), .IN4(n5966), .Q(n1246)
         );
  OA22X1 U1376 ( .IN1(n5709), .IN2(n6160), .IN3(n5719), .IN4(n1248), .Q(n1247)
         );
  OA22X1 U1377 ( .IN1(n5706), .IN2(n1249), .IN3(n5699), .IN4(n5951), .Q(n1248)
         );
  AOI22X1 U1378 ( .IN1(n5695), .IN2(\decodedPacket[2][100] ), .IN3(n5685), 
        .IN4(\decodedPacket[1][100] ), .QN(n1249) );
  OAI22X1 U1379 ( .IN1(n5767), .IN2(n6375), .IN3(n5764), .IN4(n1250), .QN(
        N9900) );
  OA22X1 U1380 ( .IN1(n5742), .IN2(n6307), .IN3(n5758), .IN4(n1251), .Q(n1250)
         );
  OA22X1 U1381 ( .IN1(n5738), .IN2(n1252), .IN3(n5730), .IN4(n6221), .Q(n1251)
         );
  OA22X1 U1382 ( .IN1(n5709), .IN2(n6153), .IN3(n5719), .IN4(n1253), .Q(n1252)
         );
  OA22X1 U1383 ( .IN1(n5706), .IN2(n1254), .IN3(n5699), .IN4(n6067), .Q(n1253)
         );
  AOI22X1 U1384 ( .IN1(n5695), .IN2(\decodedPacket[2][99] ), .IN3(n5686), 
        .IN4(\decodedPacket[1][99] ), .QN(n1254) );
  OAI22X1 U1385 ( .IN1(n5768), .IN2(n6372), .IN3(n5764), .IN4(n1255), .QN(
        N9898) );
  OA22X1 U1386 ( .IN1(n5742), .IN2(n6306), .IN3(n5759), .IN4(n1256), .Q(n1255)
         );
  OA22X1 U1387 ( .IN1(n5738), .IN2(n1257), .IN3(n5730), .IN4(n6218), .Q(n1256)
         );
  OA22X1 U1388 ( .IN1(n5709), .IN2(n6152), .IN3(n5719), .IN4(n1258), .Q(n1257)
         );
  OA22X1 U1389 ( .IN1(n5706), .IN2(n1259), .IN3(n5699), .IN4(n6064), .Q(n1258)
         );
  AOI22X1 U1390 ( .IN1(n5695), .IN2(\decodedPacket[2][98] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][98] ), .QN(n1259) );
  OAI22X1 U1391 ( .IN1(n5768), .IN2(n6377), .IN3(n5764), .IN4(n1260), .QN(
        N9896) );
  OA22X1 U1392 ( .IN1(n5741), .IN2(n6422), .IN3(n5760), .IN4(n1261), .Q(n1260)
         );
  OA22X1 U1393 ( .IN1(n5738), .IN2(n1262), .IN3(n5730), .IN4(n6223), .Q(n1261)
         );
  OA22X1 U1394 ( .IN1(n5708), .IN2(n6268), .IN3(n5719), .IN4(n1263), .Q(n1262)
         );
  OA22X1 U1395 ( .IN1(n5706), .IN2(n1264), .IN3(n5699), .IN4(n6069), .Q(n1263)
         );
  AOI22X1 U1396 ( .IN1(n5695), .IN2(\decodedPacket[2][97] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][97] ), .QN(n1264) );
  OAI22X1 U1397 ( .IN1(n5768), .IN2(n6378), .IN3(n5764), .IN4(n1265), .QN(
        N9895) );
  OA22X1 U1398 ( .IN1(n5742), .IN2(n6421), .IN3(n5756), .IN4(n1266), .Q(n1265)
         );
  OA22X1 U1399 ( .IN1(n5738), .IN2(n1267), .IN3(n5730), .IN4(n6224), .Q(n1266)
         );
  OA22X1 U1400 ( .IN1(n5709), .IN2(n6267), .IN3(n5719), .IN4(n1268), .Q(n1267)
         );
  OA22X1 U1401 ( .IN1(n5706), .IN2(n1269), .IN3(n5699), .IN4(n6070), .Q(n1268)
         );
  AOI22X1 U1402 ( .IN1(n5695), .IN2(\decodedPacket[2][96] ), .IN3(n5684), 
        .IN4(\decodedPacket[1][96] ), .QN(n1269) );
  OAI22X1 U1403 ( .IN1(n5768), .IN2(n6379), .IN3(n5764), .IN4(n1270), .QN(
        N9894) );
  OA22X1 U1404 ( .IN1(n5742), .IN2(n6420), .IN3(n5753), .IN4(n1271), .Q(n1270)
         );
  OA22X1 U1405 ( .IN1(n5738), .IN2(n1272), .IN3(n5730), .IN4(n6225), .Q(n1271)
         );
  OA22X1 U1406 ( .IN1(n5709), .IN2(n6266), .IN3(n5719), .IN4(n1273), .Q(n1272)
         );
  OA22X1 U1407 ( .IN1(n5706), .IN2(n1274), .IN3(n5699), .IN4(n6071), .Q(n1273)
         );
  AOI22X1 U1408 ( .IN1(n5695), .IN2(\decodedPacket[2][95] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][95] ), .QN(n1274) );
  OAI22X1 U1409 ( .IN1(n5768), .IN2(n6380), .IN3(n5764), .IN4(n1275), .QN(
        N9893) );
  OA22X1 U1410 ( .IN1(n5743), .IN2(n6419), .IN3(n5758), .IN4(n1276), .Q(n1275)
         );
  OA22X1 U1411 ( .IN1(n5738), .IN2(n1277), .IN3(n5730), .IN4(n6226), .Q(n1276)
         );
  OA22X1 U1412 ( .IN1(n5710), .IN2(n6265), .IN3(n5717), .IN4(n1278), .Q(n1277)
         );
  OA22X1 U1413 ( .IN1(n5706), .IN2(n1279), .IN3(n5699), .IN4(n6072), .Q(n1278)
         );
  AOI22X1 U1414 ( .IN1(n5695), .IN2(\decodedPacket[2][94] ), .IN3(n5685), 
        .IN4(\decodedPacket[1][94] ), .QN(n1279) );
  OAI22X1 U1415 ( .IN1(n5768), .IN2(n6381), .IN3(n5764), .IN4(n1280), .QN(
        N9892) );
  OA22X1 U1416 ( .IN1(n5743), .IN2(n6418), .IN3(n5758), .IN4(n1281), .Q(n1280)
         );
  OA22X1 U1417 ( .IN1(n5738), .IN2(n1282), .IN3(n5730), .IN4(n6227), .Q(n1281)
         );
  OA22X1 U1418 ( .IN1(n5710), .IN2(n6264), .IN3(n5717), .IN4(n1283), .Q(n1282)
         );
  OA22X1 U1419 ( .IN1(n5706), .IN2(n1284), .IN3(n5699), .IN4(n6073), .Q(n1283)
         );
  AOI22X1 U1420 ( .IN1(n5695), .IN2(\decodedPacket[2][93] ), .IN3(n5683), 
        .IN4(\decodedPacket[1][93] ), .QN(n1284) );
  OAI22X1 U1421 ( .IN1(n5768), .IN2(n6382), .IN3(n5764), .IN4(n1285), .QN(
        N9891) );
  OA22X1 U1422 ( .IN1(n5743), .IN2(n6417), .IN3(n5759), .IN4(n1286), .Q(n1285)
         );
  OA22X1 U1423 ( .IN1(n5738), .IN2(n1287), .IN3(n5730), .IN4(n6228), .Q(n1286)
         );
  OA22X1 U1424 ( .IN1(n5710), .IN2(n6263), .IN3(n5718), .IN4(n1288), .Q(n1287)
         );
  OA22X1 U1425 ( .IN1(n5706), .IN2(n1289), .IN3(n5699), .IN4(n6074), .Q(n1288)
         );
  AOI22X1 U1426 ( .IN1(n5695), .IN2(\decodedPacket[2][92] ), .IN3(n5685), 
        .IN4(\decodedPacket[1][92] ), .QN(n1289) );
  OAI22X1 U1427 ( .IN1(n5768), .IN2(n6383), .IN3(n5764), .IN4(n1290), .QN(
        N9890) );
  OA22X1 U1428 ( .IN1(n5743), .IN2(n6416), .IN3(n5760), .IN4(n1291), .Q(n1290)
         );
  OA22X1 U1429 ( .IN1(n5737), .IN2(n1292), .IN3(n5730), .IN4(n6229), .Q(n1291)
         );
  OA22X1 U1430 ( .IN1(n5710), .IN2(n6262), .IN3(n5720), .IN4(n1293), .Q(n1292)
         );
  OA22X1 U1431 ( .IN1(n5706), .IN2(n1294), .IN3(n5699), .IN4(n6075), .Q(n1293)
         );
  AOI22X1 U1432 ( .IN1(n5695), .IN2(\decodedPacket[2][91] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][91] ), .QN(n1294) );
  OAI22X1 U1433 ( .IN1(n5768), .IN2(n6385), .IN3(n5764), .IN4(n1295), .QN(
        N9889) );
  OA22X1 U1434 ( .IN1(n5743), .IN2(n6359), .IN3(n5756), .IN4(n1296), .Q(n1295)
         );
  OA22X1 U1435 ( .IN1(n5737), .IN2(n1297), .IN3(n5730), .IN4(n6231), .Q(n1296)
         );
  OA22X1 U1436 ( .IN1(n5710), .IN2(n6205), .IN3(n4910), .IN4(n1298), .Q(n1297)
         );
  OA22X1 U1437 ( .IN1(n5705), .IN2(n1299), .IN3(n5699), .IN4(n6077), .Q(n1298)
         );
  AOI22X1 U1438 ( .IN1(n5695), .IN2(\decodedPacket[2][90] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][90] ), .QN(n1299) );
  OAI22X1 U1439 ( .IN1(n5768), .IN2(n6386), .IN3(n5764), .IN4(n1300), .QN(
        N9888) );
  OA22X1 U1440 ( .IN1(n5743), .IN2(n6358), .IN3(n5757), .IN4(n1301), .Q(n1300)
         );
  OA22X1 U1441 ( .IN1(n5737), .IN2(n1302), .IN3(n5730), .IN4(n6232), .Q(n1301)
         );
  OA22X1 U1442 ( .IN1(n5710), .IN2(n6204), .IN3(n5724), .IN4(n1303), .Q(n1302)
         );
  OA22X1 U1443 ( .IN1(n5705), .IN2(n1304), .IN3(n5699), .IN4(n6078), .Q(n1303)
         );
  AOI22X1 U1444 ( .IN1(n5695), .IN2(\decodedPacket[2][89] ), .IN3(n5684), 
        .IN4(\decodedPacket[1][89] ), .QN(n1304) );
  OAI22X1 U1445 ( .IN1(n5768), .IN2(n6387), .IN3(n5764), .IN4(n1305), .QN(
        N9887) );
  OA22X1 U1446 ( .IN1(n5743), .IN2(n6357), .IN3(n5753), .IN4(n1306), .Q(n1305)
         );
  OA22X1 U1447 ( .IN1(n5737), .IN2(n1307), .IN3(n5730), .IN4(n6233), .Q(n1306)
         );
  OA22X1 U1448 ( .IN1(n5710), .IN2(n6203), .IN3(n5725), .IN4(n1308), .Q(n1307)
         );
  OA22X1 U1449 ( .IN1(n5705), .IN2(n1309), .IN3(n5699), .IN4(n6079), .Q(n1308)
         );
  AOI22X1 U1450 ( .IN1(n5695), .IN2(\decodedPacket[2][88] ), .IN3(n5689), 
        .IN4(\decodedPacket[1][88] ), .QN(n1309) );
  OAI22X1 U1451 ( .IN1(n5768), .IN2(n6388), .IN3(n5764), .IN4(n1310), .QN(
        N9886) );
  OA22X1 U1452 ( .IN1(n5743), .IN2(n6356), .IN3(n5754), .IN4(n1311), .Q(n1310)
         );
  OA22X1 U1453 ( .IN1(n5737), .IN2(n1312), .IN3(n5730), .IN4(n6234), .Q(n1311)
         );
  OA22X1 U1454 ( .IN1(n5710), .IN2(n6202), .IN3(n5720), .IN4(n1313), .Q(n1312)
         );
  OA22X1 U1455 ( .IN1(n5705), .IN2(n1314), .IN3(n5699), .IN4(n6080), .Q(n1313)
         );
  AOI22X1 U1456 ( .IN1(n5695), .IN2(\decodedPacket[2][87] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][87] ), .QN(n1314) );
  OAI22X1 U1457 ( .IN1(n5768), .IN2(n6389), .IN3(n5764), .IN4(n1315), .QN(
        N9885) );
  OA22X1 U1458 ( .IN1(n5742), .IN2(n6355), .IN3(n5755), .IN4(n1316), .Q(n1315)
         );
  OA22X1 U1459 ( .IN1(n5737), .IN2(n1317), .IN3(n5730), .IN4(n6235), .Q(n1316)
         );
  OA22X1 U1460 ( .IN1(n5709), .IN2(n6201), .IN3(n5723), .IN4(n1318), .Q(n1317)
         );
  OA22X1 U1461 ( .IN1(n5705), .IN2(n1319), .IN3(n5699), .IN4(n6081), .Q(n1318)
         );
  AOI22X1 U1462 ( .IN1(n5695), .IN2(\decodedPacket[2][86] ), .IN3(n5683), 
        .IN4(\decodedPacket[1][86] ), .QN(n1319) );
  OAI22X1 U1463 ( .IN1(n5769), .IN2(n6390), .IN3(n5764), .IN4(n1320), .QN(
        N9884) );
  OA22X1 U1464 ( .IN1(n5743), .IN2(n6354), .IN3(n5754), .IN4(n1321), .Q(n1320)
         );
  OA22X1 U1465 ( .IN1(n5737), .IN2(n1322), .IN3(n5730), .IN4(n6236), .Q(n1321)
         );
  OA22X1 U1466 ( .IN1(n5710), .IN2(n6200), .IN3(n5720), .IN4(n1323), .Q(n1322)
         );
  OA22X1 U1467 ( .IN1(n5705), .IN2(n1324), .IN3(n5699), .IN4(n6082), .Q(n1323)
         );
  AOI22X1 U1468 ( .IN1(n5695), .IN2(\decodedPacket[2][85] ), .IN3(n5690), 
        .IN4(\decodedPacket[1][85] ), .QN(n1324) );
  OAI22X1 U1469 ( .IN1(n5769), .IN2(n6391), .IN3(n5764), .IN4(n1325), .QN(
        N9883) );
  OA22X1 U1470 ( .IN1(n5743), .IN2(n6353), .IN3(n5755), .IN4(n1326), .Q(n1325)
         );
  OA22X1 U1471 ( .IN1(n5737), .IN2(n1327), .IN3(n5730), .IN4(n6237), .Q(n1326)
         );
  OA22X1 U1472 ( .IN1(n5710), .IN2(n6199), .IN3(n5719), .IN4(n1328), .Q(n1327)
         );
  OA22X1 U1473 ( .IN1(n5705), .IN2(n1329), .IN3(n5699), .IN4(n6083), .Q(n1328)
         );
  AOI22X1 U1474 ( .IN1(n5695), .IN2(\decodedPacket[2][84] ), .IN3(n5684), 
        .IN4(\decodedPacket[1][84] ), .QN(n1329) );
  OAI22X1 U1475 ( .IN1(n5769), .IN2(n6400), .IN3(n5764), .IN4(n1330), .QN(
        N9882) );
  OA22X1 U1476 ( .IN1(n5743), .IN2(n6415), .IN3(n5750), .IN4(n1331), .Q(n1330)
         );
  OA22X1 U1477 ( .IN1(n5737), .IN2(n1332), .IN3(n5730), .IN4(n6246), .Q(n1331)
         );
  OA22X1 U1478 ( .IN1(n5710), .IN2(n6261), .IN3(n5717), .IN4(n1333), .Q(n1332)
         );
  OA22X1 U1479 ( .IN1(n5705), .IN2(n1334), .IN3(n5699), .IN4(n6092), .Q(n1333)
         );
  AOI22X1 U1480 ( .IN1(n5694), .IN2(\decodedPacket[2][83] ), .IN3(n5686), 
        .IN4(\decodedPacket[1][83] ), .QN(n1334) );
  OAI22X1 U1481 ( .IN1(n5769), .IN2(n6406), .IN3(n5764), .IN4(n1335), .QN(
        N9881) );
  OA22X1 U1482 ( .IN1(n5743), .IN2(n6414), .IN3(n5751), .IN4(n1336), .Q(n1335)
         );
  OA22X1 U1483 ( .IN1(n5737), .IN2(n1337), .IN3(n5730), .IN4(n6252), .Q(n1336)
         );
  OA22X1 U1484 ( .IN1(n5710), .IN2(n6260), .IN3(n5726), .IN4(n1338), .Q(n1337)
         );
  OA22X1 U1485 ( .IN1(n5705), .IN2(n1339), .IN3(n5699), .IN4(n6098), .Q(n1338)
         );
  AOI22X1 U1486 ( .IN1(n5694), .IN2(\decodedPacket[2][82] ), .IN3(n5688), 
        .IN4(\decodedPacket[1][82] ), .QN(n1339) );
  OAI22X1 U1487 ( .IN1(n5769), .IN2(n6407), .IN3(n5764), .IN4(n1340), .QN(
        N9880) );
  OA22X1 U1488 ( .IN1(n5744), .IN2(n6413), .IN3(n5752), .IN4(n1341), .Q(n1340)
         );
  OA22X1 U1489 ( .IN1(n5737), .IN2(n1342), .IN3(n5730), .IN4(n6253), .Q(n1341)
         );
  OA22X1 U1490 ( .IN1(n5711), .IN2(n6259), .IN3(n5725), .IN4(n1343), .Q(n1342)
         );
  OA22X1 U1491 ( .IN1(n5705), .IN2(n1344), .IN3(n5699), .IN4(n6099), .Q(n1343)
         );
  AOI22X1 U1492 ( .IN1(n5694), .IN2(\decodedPacket[2][81] ), .IN3(n5683), 
        .IN4(\decodedPacket[1][81] ), .QN(n1344) );
  OAI22X1 U1493 ( .IN1(n5769), .IN2(n6408), .IN3(n5764), .IN4(n1345), .QN(
        N9879) );
  OA22X1 U1494 ( .IN1(n5744), .IN2(n6412), .IN3(n5757), .IN4(n1346), .Q(n1345)
         );
  OA22X1 U1495 ( .IN1(n5737), .IN2(n1347), .IN3(n5730), .IN4(n6254), .Q(n1346)
         );
  OA22X1 U1496 ( .IN1(n5711), .IN2(n6258), .IN3(n5722), .IN4(n1348), .Q(n1347)
         );
  OA22X1 U1497 ( .IN1(n5705), .IN2(n1349), .IN3(n5699), .IN4(n6100), .Q(n1348)
         );
  AOI22X1 U1498 ( .IN1(n5694), .IN2(\decodedPacket[2][80] ), .IN3(n5685), 
        .IN4(\decodedPacket[1][80] ), .QN(n1349) );
  OAI22X1 U1499 ( .IN1(n5769), .IN2(n6409), .IN3(n5764), .IN4(n1350), .QN(
        N9878) );
  OA22X1 U1500 ( .IN1(n5744), .IN2(n6411), .IN3(n5751), .IN4(n1351), .Q(n1350)
         );
  OA22X1 U1501 ( .IN1(n5736), .IN2(n1352), .IN3(n5730), .IN4(n6255), .Q(n1351)
         );
  OA22X1 U1502 ( .IN1(n5711), .IN2(n6257), .IN3(n5723), .IN4(n1353), .Q(n1352)
         );
  OA22X1 U1503 ( .IN1(n5705), .IN2(n1354), .IN3(n5699), .IN4(n6101), .Q(n1353)
         );
  AOI22X1 U1504 ( .IN1(n5694), .IN2(\decodedPacket[2][79] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][79] ), .QN(n1354) );
  OAI22X1 U1505 ( .IN1(n5769), .IN2(n6401), .IN3(n5764), .IN4(n1355), .QN(
        N9877) );
  OA22X1 U1506 ( .IN1(n5744), .IN2(n6410), .IN3(n5753), .IN4(n1356), .Q(n1355)
         );
  OA22X1 U1507 ( .IN1(n5736), .IN2(n1357), .IN3(n5731), .IN4(n6247), .Q(n1356)
         );
  OA22X1 U1508 ( .IN1(n5711), .IN2(n6256), .IN3(n5726), .IN4(n1358), .Q(n1357)
         );
  OA22X1 U1509 ( .IN1(n5705), .IN2(n1359), .IN3(n5699), .IN4(n6093), .Q(n1358)
         );
  AOI22X1 U1510 ( .IN1(n5694), .IN2(\decodedPacket[2][78] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][78] ), .QN(n1359) );
  OAI22X1 U1511 ( .IN1(n5769), .IN2(n6399), .IN3(n5764), .IN4(n1360), .QN(
        N9876) );
  OA22X1 U1512 ( .IN1(n5744), .IN2(n6352), .IN3(n5756), .IN4(n1361), .Q(n1360)
         );
  OA22X1 U1513 ( .IN1(n5736), .IN2(n1362), .IN3(n5731), .IN4(n6244), .Q(n1361)
         );
  OA22X1 U1514 ( .IN1(n5711), .IN2(n6198), .IN3(n5724), .IN4(n1363), .Q(n1362)
         );
  OA22X1 U1515 ( .IN1(n5705), .IN2(n1364), .IN3(n5700), .IN4(n6090), .Q(n1363)
         );
  AOI22X1 U1516 ( .IN1(n5694), .IN2(\decodedPacket[2][77] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][77] ), .QN(n1364) );
  OAI22X1 U1517 ( .IN1(n5769), .IN2(n6398), .IN3(n5764), .IN4(n1365), .QN(
        N9875) );
  OA22X1 U1518 ( .IN1(n5744), .IN2(n6402), .IN3(n5750), .IN4(n1366), .Q(n1365)
         );
  OA22X1 U1519 ( .IN1(n5736), .IN2(n1367), .IN3(n5731), .IN4(n6243), .Q(n1366)
         );
  OA22X1 U1520 ( .IN1(n5711), .IN2(n6248), .IN3(n5721), .IN4(n1368), .Q(n1367)
         );
  OA22X1 U1521 ( .IN1(n5704), .IN2(n1369), .IN3(n5700), .IN4(n6089), .Q(n1368)
         );
  AOI22X1 U1522 ( .IN1(n5694), .IN2(\decodedPacket[2][76] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][76] ), .QN(n1369) );
  OAI22X1 U1523 ( .IN1(n5769), .IN2(n6397), .IN3(n5764), .IN4(n1370), .QN(
        N9874) );
  OA22X1 U1524 ( .IN1(n5744), .IN2(n6403), .IN3(n5752), .IN4(n1371), .Q(n1370)
         );
  OA22X1 U1525 ( .IN1(n5736), .IN2(n1372), .IN3(n5731), .IN4(n6242), .Q(n1371)
         );
  OA22X1 U1526 ( .IN1(n5711), .IN2(n6249), .IN3(n5720), .IN4(n1373), .Q(n1372)
         );
  OA22X1 U1527 ( .IN1(n5704), .IN2(n1374), .IN3(n5700), .IN4(n6087), .Q(n1373)
         );
  AOI22X1 U1528 ( .IN1(n5694), .IN2(\decodedPacket[2][75] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][75] ), .QN(n1374) );
  OAI22X1 U1529 ( .IN1(n5769), .IN2(n6396), .IN3(n5765), .IN4(n1375), .QN(
        N9873) );
  OA22X1 U1530 ( .IN1(n5743), .IN2(n6404), .IN3(n5754), .IN4(n1376), .Q(n1375)
         );
  OA22X1 U1531 ( .IN1(n5736), .IN2(n1377), .IN3(n5731), .IN4(n6241), .Q(n1376)
         );
  OA22X1 U1532 ( .IN1(n5710), .IN2(n6250), .IN3(n4910), .IN4(n1378), .Q(n1377)
         );
  OA22X1 U1533 ( .IN1(n5704), .IN2(n1379), .IN3(n5700), .IN4(n6088), .Q(n1378)
         );
  AOI22X1 U1534 ( .IN1(n5694), .IN2(\decodedPacket[2][74] ), .IN3(n5687), 
        .IN4(\decodedPacket[1][74] ), .QN(n1379) );
  OAI22X1 U1535 ( .IN1(n5770), .IN2(n6396), .IN3(n5765), .IN4(n1380), .QN(
        N9872) );
  OA22X1 U1536 ( .IN1(n5744), .IN2(n6405), .IN3(n5751), .IN4(n1381), .Q(n1380)
         );
  OA22X1 U1537 ( .IN1(n5736), .IN2(n1382), .IN3(n5731), .IN4(n6242), .Q(n1381)
         );
  OA22X1 U1538 ( .IN1(n5711), .IN2(n6251), .IN3(n5718), .IN4(n1383), .Q(n1382)
         );
  OA22X1 U1539 ( .IN1(n5704), .IN2(n1384), .IN3(n5700), .IN4(n6087), .Q(n1383)
         );
  AOI22X1 U1540 ( .IN1(n5694), .IN2(\decodedPacket[2][73] ), .IN3(n5686), 
        .IN4(\decodedPacket[1][73] ), .QN(n1384) );
  OAI22X1 U1541 ( .IN1(n5769), .IN2(n6394), .IN3(n5765), .IN4(n1385), .QN(
        N9871) );
  OA22X1 U1542 ( .IN1(n5744), .IN2(n6393), .IN3(n5760), .IN4(n1386), .Q(n1385)
         );
  OA22X1 U1543 ( .IN1(n5736), .IN2(n1387), .IN3(n5731), .IN4(n6240), .Q(n1386)
         );
  OA22X1 U1544 ( .IN1(n5711), .IN2(n6239), .IN3(n5717), .IN4(n1388), .Q(n1387)
         );
  OA22X1 U1545 ( .IN1(n5704), .IN2(n1389), .IN3(n5700), .IN4(n6086), .Q(n1388)
         );
  AOI22X1 U1546 ( .IN1(n5694), .IN2(\decodedPacket[2][72] ), .IN3(n5686), 
        .IN4(\decodedPacket[1][72] ), .QN(n1389) );
  OAI22X1 U1547 ( .IN1(n5770), .IN2(n6361), .IN3(n5765), .IN4(n1390), .QN(
        N9870) );
  OA22X1 U1548 ( .IN1(n5744), .IN2(n6360), .IN3(n5756), .IN4(n1391), .Q(n1390)
         );
  OA22X1 U1549 ( .IN1(n5736), .IN2(n1392), .IN3(n5731), .IN4(n6207), .Q(n1391)
         );
  OA22X1 U1550 ( .IN1(n5711), .IN2(n6206), .IN3(n5718), .IN4(n1393), .Q(n1392)
         );
  OA22X1 U1551 ( .IN1(n5704), .IN2(n1394), .IN3(n5700), .IN4(n6053), .Q(n1393)
         );
  AOI22X1 U1552 ( .IN1(n5694), .IN2(\decodedPacket[2][71] ), .IN3(n5686), 
        .IN4(\decodedPacket[1][71] ), .QN(n1394) );
  OAI22X1 U1553 ( .IN1(n6350), .IN2(n5770), .IN3(n5765), .IN4(n1395), .QN(
        N9869) );
  OA22X1 U1554 ( .IN1(n6351), .IN2(n5744), .IN3(n5756), .IN4(n1396), .Q(n1395)
         );
  OA22X1 U1555 ( .IN1(n5736), .IN2(n1397), .IN3(n6196), .IN4(n5731), .Q(n1396)
         );
  OA22X1 U1556 ( .IN1(n6197), .IN2(n5711), .IN3(n5726), .IN4(n1398), .Q(n1397)
         );
  OA22X1 U1557 ( .IN1(n5704), .IN2(n1399), .IN3(n6042), .IN4(n5700), .Q(n1398)
         );
  AOI22X1 U1558 ( .IN1(\decodedPacket[2][70] ), .IN2(n5694), .IN3(n5686), 
        .IN4(\decodedPacket[1][70] ), .QN(n1399) );
  OAI22X1 U1559 ( .IN1(n6395), .IN2(n5770), .IN3(n5765), .IN4(n1400), .QN(
        N9868) );
  OA22X1 U1560 ( .IN1(n6392), .IN2(n5744), .IN3(n5757), .IN4(n1401), .Q(n1400)
         );
  OA22X1 U1561 ( .IN1(n5736), .IN2(n1402), .IN3(n6242), .IN4(n5731), .Q(n1401)
         );
  OA22X1 U1562 ( .IN1(n6238), .IN2(n5711), .IN3(n5726), .IN4(n1403), .Q(n1402)
         );
  OA22X1 U1563 ( .IN1(n5704), .IN2(n1404), .IN3(n6088), .IN4(n5700), .Q(n1403)
         );
  AOI22X1 U1564 ( .IN1(\decodedPacket[2][69] ), .IN2(n5694), .IN3(n5686), 
        .IN4(\decodedPacket[1][69] ), .QN(n1404) );
  OAI22X1 U1565 ( .IN1(n6423), .IN2(n5770), .IN3(n5765), .IN4(n1405), .QN(
        N9867) );
  OA22X1 U1566 ( .IN1(n6423), .IN2(n5744), .IN3(n5758), .IN4(n1406), .Q(n1405)
         );
  OA22X1 U1567 ( .IN1(n5736), .IN2(n1407), .IN3(n6269), .IN4(n5731), .Q(n1406)
         );
  OA22X1 U1568 ( .IN1(n6269), .IN2(n5711), .IN3(n5717), .IN4(n1408), .Q(n1407)
         );
  OA22X1 U1569 ( .IN1(n5704), .IN2(n1409), .IN3(n6115), .IN4(n5700), .Q(n1408)
         );
  AOI22X1 U1570 ( .IN1(\decodedPacket[2][68] ), .IN2(n5694), .IN3(n5686), 
        .IN4(\decodedPacket[1][68] ), .QN(n1409) );
  OAI22X1 U1571 ( .IN1(n6424), .IN2(n5770), .IN3(n5765), .IN4(n1410), .QN(
        N9866) );
  OA22X1 U1572 ( .IN1(n6424), .IN2(n5745), .IN3(n5753), .IN4(n1411), .Q(n1410)
         );
  OA22X1 U1573 ( .IN1(n5735), .IN2(n1412), .IN3(n6270), .IN4(n5731), .Q(n1411)
         );
  OA22X1 U1574 ( .IN1(n6270), .IN2(n5712), .IN3(n5718), .IN4(n1413), .Q(n1412)
         );
  OA22X1 U1575 ( .IN1(n5704), .IN2(n1414), .IN3(n6116), .IN4(n5700), .Q(n1413)
         );
  AOI22X1 U1576 ( .IN1(\decodedPacket[2][67] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][67] ), .QN(n1414) );
  OAI22X1 U1577 ( .IN1(n6425), .IN2(n5770), .IN3(n5765), .IN4(n1415), .QN(
        N9865) );
  OA22X1 U1578 ( .IN1(n6425), .IN2(n5745), .IN3(n5758), .IN4(n1416), .Q(n1415)
         );
  OA22X1 U1579 ( .IN1(n5735), .IN2(n1417), .IN3(n6271), .IN4(n5731), .Q(n1416)
         );
  OA22X1 U1580 ( .IN1(n6271), .IN2(n5712), .IN3(n5721), .IN4(n1418), .Q(n1417)
         );
  OA22X1 U1581 ( .IN1(n5704), .IN2(n1419), .IN3(n6117), .IN4(n5700), .Q(n1418)
         );
  AOI22X1 U1582 ( .IN1(\decodedPacket[2][66] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][66] ), .QN(n1419) );
  OAI22X1 U1583 ( .IN1(n6426), .IN2(n5770), .IN3(n5765), .IN4(n1420), .QN(
        N9864) );
  OA22X1 U1584 ( .IN1(n6426), .IN2(n5745), .IN3(n5753), .IN4(n1421), .Q(n1420)
         );
  OA22X1 U1585 ( .IN1(n5735), .IN2(n1422), .IN3(n6272), .IN4(n5731), .Q(n1421)
         );
  OA22X1 U1586 ( .IN1(n6272), .IN2(n5712), .IN3(n5720), .IN4(n1423), .Q(n1422)
         );
  OA22X1 U1587 ( .IN1(n5704), .IN2(n1424), .IN3(n6118), .IN4(n5700), .Q(n1423)
         );
  AOI22X1 U1588 ( .IN1(\decodedPacket[2][65] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][65] ), .QN(n1424) );
  OAI22X1 U1589 ( .IN1(n6427), .IN2(n5770), .IN3(n5765), .IN4(n1425), .QN(
        N9863) );
  OA22X1 U1590 ( .IN1(n6427), .IN2(n5745), .IN3(n5759), .IN4(n1426), .Q(n1425)
         );
  OA22X1 U1591 ( .IN1(n5735), .IN2(n1427), .IN3(n6273), .IN4(n5731), .Q(n1426)
         );
  OA22X1 U1592 ( .IN1(n6273), .IN2(n5712), .IN3(n5723), .IN4(n1428), .Q(n1427)
         );
  OA22X1 U1593 ( .IN1(n5704), .IN2(n1429), .IN3(n6119), .IN4(n5700), .Q(n1428)
         );
  AOI22X1 U1594 ( .IN1(\decodedPacket[2][64] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][64] ), .QN(n1429) );
  OAI22X1 U1595 ( .IN1(n6428), .IN2(n5770), .IN3(n5765), .IN4(n1430), .QN(
        N9862) );
  OA22X1 U1596 ( .IN1(n6428), .IN2(n5745), .IN3(n5758), .IN4(n1431), .Q(n1430)
         );
  OA22X1 U1597 ( .IN1(n5735), .IN2(n1432), .IN3(n6274), .IN4(n5731), .Q(n1431)
         );
  OA22X1 U1598 ( .IN1(n6274), .IN2(n5712), .IN3(n5725), .IN4(n1433), .Q(n1432)
         );
  OA22X1 U1599 ( .IN1(n5704), .IN2(n1434), .IN3(n6120), .IN4(n5700), .Q(n1433)
         );
  AOI22X1 U1600 ( .IN1(\decodedPacket[2][63] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][63] ), .QN(n1434) );
  OAI22X1 U1601 ( .IN1(n6429), .IN2(n5770), .IN3(n5765), .IN4(n1435), .QN(
        N9861) );
  OA22X1 U1602 ( .IN1(n6429), .IN2(n5745), .IN3(n5760), .IN4(n1436), .Q(n1435)
         );
  OA22X1 U1603 ( .IN1(n5735), .IN2(n1437), .IN3(n6275), .IN4(n5731), .Q(n1436)
         );
  OA22X1 U1604 ( .IN1(n6275), .IN2(n5712), .IN3(n5719), .IN4(n1438), .Q(n1437)
         );
  OA22X1 U1605 ( .IN1(n5704), .IN2(n1439), .IN3(n6121), .IN4(n5700), .Q(n1438)
         );
  AOI22X1 U1606 ( .IN1(\decodedPacket[2][62] ), .IN2(n5694), .IN3(n5685), 
        .IN4(\decodedPacket[1][62] ), .QN(n1439) );
  OAI22X1 U1607 ( .IN1(n6430), .IN2(n5770), .IN3(n5765), .IN4(n1440), .QN(
        N9860) );
  OA22X1 U1608 ( .IN1(n6430), .IN2(n5745), .IN3(n5755), .IN4(n1441), .Q(n1440)
         );
  OA22X1 U1609 ( .IN1(n5735), .IN2(n1442), .IN3(n6276), .IN4(n5731), .Q(n1441)
         );
  OA22X1 U1610 ( .IN1(n6276), .IN2(n5712), .IN3(n4910), .IN4(n1443), .Q(n1442)
         );
  OA22X1 U1611 ( .IN1(n5703), .IN2(n1444), .IN3(n6122), .IN4(n5700), .Q(n1443)
         );
  AOI22X1 U1612 ( .IN1(\decodedPacket[2][61] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][61] ), .QN(n1444) );
  OAI22X1 U1613 ( .IN1(n6431), .IN2(n5770), .IN3(n5765), .IN4(n1445), .QN(
        N9859) );
  OA22X1 U1614 ( .IN1(n6431), .IN2(n5745), .IN3(n5755), .IN4(n1446), .Q(n1445)
         );
  OA22X1 U1615 ( .IN1(n5735), .IN2(n1447), .IN3(n6277), .IN4(n5731), .Q(n1446)
         );
  OA22X1 U1616 ( .IN1(n6277), .IN2(n5712), .IN3(n5724), .IN4(n1448), .Q(n1447)
         );
  OA22X1 U1617 ( .IN1(n5703), .IN2(n1449), .IN3(n6123), .IN4(n5700), .Q(n1448)
         );
  AOI22X1 U1618 ( .IN1(\decodedPacket[2][60] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][60] ), .QN(n1449) );
  OAI22X1 U1619 ( .IN1(n6432), .IN2(n5770), .IN3(n5765), .IN4(n1450), .QN(
        N9858) );
  OA22X1 U1620 ( .IN1(n6432), .IN2(n5745), .IN3(n5752), .IN4(n1451), .Q(n1450)
         );
  OA22X1 U1621 ( .IN1(n5735), .IN2(n1452), .IN3(n6278), .IN4(n5731), .Q(n1451)
         );
  OA22X1 U1622 ( .IN1(n6278), .IN2(n5712), .IN3(n5722), .IN4(n1453), .Q(n1452)
         );
  OA22X1 U1623 ( .IN1(n5703), .IN2(n1454), .IN3(n6124), .IN4(n5700), .Q(n1453)
         );
  AOI22X1 U1624 ( .IN1(\decodedPacket[2][59] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][59] ), .QN(n1454) );
  OAI22X1 U1625 ( .IN1(n6433), .IN2(n5771), .IN3(n5765), .IN4(n1455), .QN(
        N9857) );
  OA22X1 U1626 ( .IN1(n6433), .IN2(n5745), .IN3(n5754), .IN4(n1456), .Q(n1455)
         );
  OA22X1 U1627 ( .IN1(n5735), .IN2(n1457), .IN3(n6279), .IN4(n5731), .Q(n1456)
         );
  OA22X1 U1628 ( .IN1(n6279), .IN2(n5712), .IN3(n5717), .IN4(n1458), .Q(n1457)
         );
  OA22X1 U1629 ( .IN1(n5703), .IN2(n1459), .IN3(n6125), .IN4(n5700), .Q(n1458)
         );
  AOI22X1 U1630 ( .IN1(\decodedPacket[2][58] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][58] ), .QN(n1459) );
  OAI22X1 U1631 ( .IN1(n6434), .IN2(n5771), .IN3(n5765), .IN4(n1460), .QN(
        N9856) );
  OA22X1 U1632 ( .IN1(n6434), .IN2(n5745), .IN3(n5750), .IN4(n1461), .Q(n1460)
         );
  OA22X1 U1633 ( .IN1(n5735), .IN2(n1462), .IN3(n6280), .IN4(n5731), .Q(n1461)
         );
  OA22X1 U1634 ( .IN1(n6280), .IN2(n5712), .IN3(n5718), .IN4(n1463), .Q(n1462)
         );
  OA22X1 U1635 ( .IN1(n5703), .IN2(n1464), .IN3(n6126), .IN4(n5700), .Q(n1463)
         );
  AOI22X1 U1636 ( .IN1(\decodedPacket[2][57] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][57] ), .QN(n1464) );
  OAI22X1 U1637 ( .IN1(n6435), .IN2(n5771), .IN3(n5765), .IN4(n1465), .QN(
        N9855) );
  OA22X1 U1638 ( .IN1(n6435), .IN2(n5745), .IN3(n5751), .IN4(n1466), .Q(n1465)
         );
  OA22X1 U1639 ( .IN1(n5735), .IN2(n1467), .IN3(n6281), .IN4(n5731), .Q(n1466)
         );
  OA22X1 U1640 ( .IN1(n6281), .IN2(n5712), .IN3(n5721), .IN4(n1468), .Q(n1467)
         );
  OA22X1 U1641 ( .IN1(n5703), .IN2(n1469), .IN3(n6127), .IN4(n5700), .Q(n1468)
         );
  AOI22X1 U1642 ( .IN1(\decodedPacket[2][56] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][56] ), .QN(n1469) );
  OAI22X1 U1643 ( .IN1(n6436), .IN2(n5771), .IN3(n5765), .IN4(n1470), .QN(
        N9854) );
  OA22X1 U1644 ( .IN1(n6436), .IN2(n5745), .IN3(n5750), .IN4(n1471), .Q(n1470)
         );
  OA22X1 U1645 ( .IN1(n5734), .IN2(n1472), .IN3(n6282), .IN4(n5731), .Q(n1471)
         );
  OA22X1 U1646 ( .IN1(n6282), .IN2(n5712), .IN3(n5722), .IN4(n1473), .Q(n1472)
         );
  OA22X1 U1647 ( .IN1(n5703), .IN2(n1474), .IN3(n6128), .IN4(n5700), .Q(n1473)
         );
  AOI22X1 U1648 ( .IN1(\decodedPacket[2][55] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][55] ), .QN(n1474) );
  OAI22X1 U1649 ( .IN1(n6437), .IN2(n5771), .IN3(n5765), .IN4(n1475), .QN(
        N9853) );
  OA22X1 U1650 ( .IN1(n6437), .IN2(n5746), .IN3(n5750), .IN4(n1476), .Q(n1475)
         );
  OA22X1 U1651 ( .IN1(n5734), .IN2(n1477), .IN3(n6283), .IN4(n5731), .Q(n1476)
         );
  OA22X1 U1652 ( .IN1(n6283), .IN2(n5713), .IN3(n5721), .IN4(n1478), .Q(n1477)
         );
  OA22X1 U1653 ( .IN1(n5703), .IN2(n1479), .IN3(n6129), .IN4(n5700), .Q(n1478)
         );
  AOI22X1 U1654 ( .IN1(\decodedPacket[2][54] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][54] ), .QN(n1479) );
  OAI22X1 U1655 ( .IN1(n6438), .IN2(n5771), .IN3(n5765), .IN4(n1480), .QN(
        N9852) );
  OA22X1 U1656 ( .IN1(n6438), .IN2(n5746), .IN3(n5750), .IN4(n1481), .Q(n1480)
         );
  OA22X1 U1657 ( .IN1(n5734), .IN2(n1482), .IN3(n6284), .IN4(n5731), .Q(n1481)
         );
  OA22X1 U1658 ( .IN1(n6284), .IN2(n5713), .IN3(n4910), .IN4(n1483), .Q(n1482)
         );
  OA22X1 U1659 ( .IN1(n5703), .IN2(n1484), .IN3(n6130), .IN4(n5700), .Q(n1483)
         );
  AOI22X1 U1660 ( .IN1(\decodedPacket[2][53] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][53] ), .QN(n1484) );
  OAI22X1 U1661 ( .IN1(n6439), .IN2(n5771), .IN3(n5765), .IN4(n1485), .QN(
        N9851) );
  OA22X1 U1662 ( .IN1(n6439), .IN2(n5746), .IN3(n5750), .IN4(n1486), .Q(n1485)
         );
  OA22X1 U1663 ( .IN1(n5734), .IN2(n1487), .IN3(n6285), .IN4(n5731), .Q(n1486)
         );
  OA22X1 U1664 ( .IN1(n6285), .IN2(n5713), .IN3(n4910), .IN4(n1488), .Q(n1487)
         );
  OA22X1 U1665 ( .IN1(n5703), .IN2(n1489), .IN3(n6131), .IN4(n5700), .Q(n1488)
         );
  AOI22X1 U1666 ( .IN1(\decodedPacket[2][52] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][52] ), .QN(n1489) );
  OAI22X1 U1667 ( .IN1(n6440), .IN2(n5771), .IN3(n5765), .IN4(n1490), .QN(
        N9850) );
  OA22X1 U1668 ( .IN1(n6440), .IN2(n5746), .IN3(n5750), .IN4(n1491), .Q(n1490)
         );
  OA22X1 U1669 ( .IN1(n5734), .IN2(n1492), .IN3(n6286), .IN4(n5731), .Q(n1491)
         );
  OA22X1 U1670 ( .IN1(n6286), .IN2(n5713), .IN3(n5724), .IN4(n1493), .Q(n1492)
         );
  OA22X1 U1671 ( .IN1(n5703), .IN2(n1494), .IN3(n6132), .IN4(n5700), .Q(n1493)
         );
  AOI22X1 U1672 ( .IN1(\decodedPacket[2][51] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][51] ), .QN(n1494) );
  OAI22X1 U1673 ( .IN1(n6441), .IN2(n5771), .IN3(n5765), .IN4(n1495), .QN(
        N9849) );
  OA22X1 U1674 ( .IN1(n6441), .IN2(n5746), .IN3(n5751), .IN4(n1496), .Q(n1495)
         );
  OA22X1 U1675 ( .IN1(n5734), .IN2(n1497), .IN3(n6287), .IN4(n5731), .Q(n1496)
         );
  OA22X1 U1676 ( .IN1(n6287), .IN2(n5713), .IN3(n5720), .IN4(n1498), .Q(n1497)
         );
  OA22X1 U1677 ( .IN1(n5703), .IN2(n1499), .IN3(n6133), .IN4(n5700), .Q(n1498)
         );
  AOI22X1 U1678 ( .IN1(\decodedPacket[2][50] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][50] ), .QN(n1499) );
  OAI22X1 U1679 ( .IN1(n6442), .IN2(n5771), .IN3(n5765), .IN4(n1500), .QN(
        N9848) );
  OA22X1 U1680 ( .IN1(n6442), .IN2(n5746), .IN3(n5751), .IN4(n1501), .Q(n1500)
         );
  OA22X1 U1681 ( .IN1(n5734), .IN2(n1502), .IN3(n6288), .IN4(n5731), .Q(n1501)
         );
  OA22X1 U1682 ( .IN1(n6288), .IN2(n5713), .IN3(n5720), .IN4(n1503), .Q(n1502)
         );
  OA22X1 U1683 ( .IN1(n5703), .IN2(n1504), .IN3(n6134), .IN4(n5700), .Q(n1503)
         );
  AOI22X1 U1684 ( .IN1(\decodedPacket[2][49] ), .IN2(n5694), .IN3(n5690), 
        .IN4(\decodedPacket[1][49] ), .QN(n1504) );
  OAI22X1 U1685 ( .IN1(n6443), .IN2(n5771), .IN3(n5765), .IN4(n1505), .QN(
        N9846) );
  OA22X1 U1686 ( .IN1(n6443), .IN2(n5746), .IN3(n5751), .IN4(n1506), .Q(n1505)
         );
  OA22X1 U1687 ( .IN1(n5734), .IN2(n1507), .IN3(n6289), .IN4(n5731), .Q(n1506)
         );
  OA22X1 U1688 ( .IN1(n6289), .IN2(n5713), .IN3(n5720), .IN4(n1508), .Q(n1507)
         );
  OA22X1 U1689 ( .IN1(n5703), .IN2(n1509), .IN3(n6135), .IN4(n5700), .Q(n1508)
         );
  AOI22X1 U1690 ( .IN1(\decodedPacket[2][48] ), .IN2(n5694), .IN3(n5690), 
        .IN4(\decodedPacket[1][48] ), .QN(n1509) );
  OAI22X1 U1691 ( .IN1(n6444), .IN2(n5771), .IN3(n5765), .IN4(n1510), .QN(
        N9845) );
  OA22X1 U1692 ( .IN1(n6444), .IN2(n5746), .IN3(n5751), .IN4(n1511), .Q(n1510)
         );
  OA22X1 U1693 ( .IN1(n5734), .IN2(n1512), .IN3(n6290), .IN4(n5731), .Q(n1511)
         );
  OA22X1 U1694 ( .IN1(n6290), .IN2(n5713), .IN3(n5720), .IN4(n1513), .Q(n1512)
         );
  OA22X1 U1695 ( .IN1(n5703), .IN2(n1514), .IN3(n6136), .IN4(n5700), .Q(n1513)
         );
  AOI22X1 U1696 ( .IN1(\decodedPacket[2][47] ), .IN2(n5694), .IN3(n5687), 
        .IN4(\decodedPacket[1][47] ), .QN(n1514) );
  OAI22X1 U1697 ( .IN1(n6445), .IN2(n5771), .IN3(n5765), .IN4(n1515), .QN(
        N9844) );
  OA22X1 U1698 ( .IN1(n6445), .IN2(n5746), .IN3(n5751), .IN4(n1516), .Q(n1515)
         );
  OA22X1 U1699 ( .IN1(n5734), .IN2(n1517), .IN3(n6291), .IN4(n5731), .Q(n1516)
         );
  OA22X1 U1700 ( .IN1(n6291), .IN2(n5713), .IN3(n5720), .IN4(n1518), .Q(n1517)
         );
  OA22X1 U1701 ( .IN1(n5702), .IN2(n1519), .IN3(n6137), .IN4(n5700), .Q(n1518)
         );
  AOI22X1 U1702 ( .IN1(\decodedPacket[2][46] ), .IN2(n5694), .IN3(n5688), 
        .IN4(\decodedPacket[1][46] ), .QN(n1519) );
  OAI22X1 U1703 ( .IN1(n6446), .IN2(n5771), .IN3(n5765), .IN4(n1520), .QN(
        N9843) );
  OA22X1 U1704 ( .IN1(n6446), .IN2(n5746), .IN3(n5752), .IN4(n1521), .Q(n1520)
         );
  OA22X1 U1705 ( .IN1(n5734), .IN2(n1522), .IN3(n6292), .IN4(n5731), .Q(n1521)
         );
  OA22X1 U1706 ( .IN1(n6292), .IN2(n5713), .IN3(n5721), .IN4(n1523), .Q(n1522)
         );
  OA22X1 U1707 ( .IN1(n5702), .IN2(n1524), .IN3(n6138), .IN4(n5700), .Q(n1523)
         );
  AOI22X1 U1708 ( .IN1(\decodedPacket[2][45] ), .IN2(n5694), .IN3(n5683), 
        .IN4(\decodedPacket[1][45] ), .QN(n1524) );
  OAI22X1 U1709 ( .IN1(n6447), .IN2(n5771), .IN3(n5765), .IN4(n1525), .QN(
        N9842) );
  OA22X1 U1710 ( .IN1(n6447), .IN2(n5746), .IN3(n5752), .IN4(n1526), .Q(n1525)
         );
  OA22X1 U1711 ( .IN1(n5734), .IN2(n1527), .IN3(n6293), .IN4(n5732), .Q(n1526)
         );
  OA22X1 U1712 ( .IN1(n6293), .IN2(n5713), .IN3(n5721), .IN4(n1528), .Q(n1527)
         );
  OA22X1 U1713 ( .IN1(n5702), .IN2(n1529), .IN3(n6139), .IN4(n5700), .Q(n1528)
         );
  AOI22X1 U1714 ( .IN1(\decodedPacket[2][44] ), .IN2(n5694), .IN3(n5684), 
        .IN4(\decodedPacket[1][44] ), .QN(n1529) );
  OAI22X1 U1715 ( .IN1(n6448), .IN2(n5771), .IN3(n5765), .IN4(n1530), .QN(
        N9841) );
  OA22X1 U1716 ( .IN1(n6448), .IN2(n5746), .IN3(n5752), .IN4(n1531), .Q(n1530)
         );
  OA22X1 U1717 ( .IN1(n5733), .IN2(n1532), .IN3(n6294), .IN4(n5732), .Q(n1531)
         );
  OA22X1 U1718 ( .IN1(n6294), .IN2(n5713), .IN3(n5721), .IN4(n1533), .Q(n1532)
         );
  OA22X1 U1719 ( .IN1(n5702), .IN2(n1534), .IN3(n6140), .IN4(n5701), .Q(n1533)
         );
  AOI22X1 U1720 ( .IN1(\decodedPacket[2][43] ), .IN2(n5694), .IN3(n5686), 
        .IN4(\decodedPacket[1][43] ), .QN(n1534) );
  OAI22X1 U1721 ( .IN1(n6449), .IN2(n5772), .IN3(n5765), .IN4(n1535), .QN(
        N9840) );
  OA22X1 U1722 ( .IN1(n6449), .IN2(n5746), .IN3(n5752), .IN4(n1536), .Q(n1535)
         );
  OA22X1 U1723 ( .IN1(n5733), .IN2(n1537), .IN3(n6295), .IN4(n5732), .Q(n1536)
         );
  OA22X1 U1724 ( .IN1(n6295), .IN2(n5713), .IN3(n5721), .IN4(n1538), .Q(n1537)
         );
  OA22X1 U1725 ( .IN1(n5702), .IN2(n1539), .IN3(n6141), .IN4(n5701), .Q(n1538)
         );
  AOI22X1 U1726 ( .IN1(\decodedPacket[2][42] ), .IN2(n5694), .IN3(n5687), 
        .IN4(\decodedPacket[1][42] ), .QN(n1539) );
  OAI22X1 U1727 ( .IN1(n6450), .IN2(n5772), .IN3(n5765), .IN4(n1540), .QN(
        N9839) );
  OA22X1 U1728 ( .IN1(n6450), .IN2(n5746), .IN3(n5752), .IN4(n1541), .Q(n1540)
         );
  OA22X1 U1729 ( .IN1(n5733), .IN2(n1542), .IN3(n6296), .IN4(n5732), .Q(n1541)
         );
  OA22X1 U1730 ( .IN1(n6296), .IN2(n5713), .IN3(n5721), .IN4(n1543), .Q(n1542)
         );
  OA22X1 U1731 ( .IN1(n5702), .IN2(n1544), .IN3(n6142), .IN4(n5701), .Q(n1543)
         );
  AOI22X1 U1732 ( .IN1(\decodedPacket[2][41] ), .IN2(n5694), .IN3(n5689), 
        .IN4(\decodedPacket[1][41] ), .QN(n1544) );
  OAI22X1 U1733 ( .IN1(n6451), .IN2(n5772), .IN3(n5765), .IN4(n1545), .QN(
        N9838) );
  OA22X1 U1734 ( .IN1(n6451), .IN2(n5747), .IN3(n5753), .IN4(n1546), .Q(n1545)
         );
  OA22X1 U1735 ( .IN1(n5733), .IN2(n1547), .IN3(n6297), .IN4(n5732), .Q(n1546)
         );
  OA22X1 U1736 ( .IN1(n6297), .IN2(n5714), .IN3(n5722), .IN4(n1548), .Q(n1547)
         );
  OA22X1 U1737 ( .IN1(n5702), .IN2(n1549), .IN3(n6143), .IN4(n5701), .Q(n1548)
         );
  AOI22X1 U1738 ( .IN1(\decodedPacket[2][40] ), .IN2(n5694), .IN3(n5687), 
        .IN4(\decodedPacket[1][40] ), .QN(n1549) );
  OAI22X1 U1739 ( .IN1(n6452), .IN2(n5772), .IN3(n5765), .IN4(n1550), .QN(
        N9837) );
  OA22X1 U1740 ( .IN1(n6452), .IN2(n5747), .IN3(n5753), .IN4(n1551), .Q(n1550)
         );
  OA22X1 U1741 ( .IN1(n5733), .IN2(n1552), .IN3(n6298), .IN4(n5732), .Q(n1551)
         );
  OA22X1 U1742 ( .IN1(n6298), .IN2(n5714), .IN3(n5722), .IN4(n1553), .Q(n1552)
         );
  OA22X1 U1743 ( .IN1(n5702), .IN2(n1554), .IN3(n6144), .IN4(n5701), .Q(n1553)
         );
  AOI22X1 U1744 ( .IN1(\decodedPacket[2][39] ), .IN2(n5694), .IN3(n5689), 
        .IN4(\decodedPacket[1][39] ), .QN(n1554) );
  OAI22X1 U1745 ( .IN1(n6453), .IN2(n5772), .IN3(n5765), .IN4(n1555), .QN(
        N9836) );
  OA22X1 U1746 ( .IN1(n6453), .IN2(n5747), .IN3(n5753), .IN4(n1556), .Q(n1555)
         );
  OA22X1 U1747 ( .IN1(n5733), .IN2(n1557), .IN3(n6299), .IN4(n5732), .Q(n1556)
         );
  OA22X1 U1748 ( .IN1(n6299), .IN2(n5714), .IN3(n5722), .IN4(n1558), .Q(n1557)
         );
  OA22X1 U1749 ( .IN1(n5702), .IN2(n1559), .IN3(n6145), .IN4(n5701), .Q(n1558)
         );
  AOI22X1 U1750 ( .IN1(\decodedPacket[2][38] ), .IN2(n5693), .IN3(n5685), 
        .IN4(\decodedPacket[1][38] ), .QN(n1559) );
  OAI22X1 U1751 ( .IN1(n6454), .IN2(n5772), .IN3(n5765), .IN4(n1560), .QN(
        N9835) );
  OA22X1 U1752 ( .IN1(n6454), .IN2(n5747), .IN3(n5753), .IN4(n1561), .Q(n1560)
         );
  OA22X1 U1753 ( .IN1(n5733), .IN2(n1562), .IN3(n6300), .IN4(n5732), .Q(n1561)
         );
  OA22X1 U1754 ( .IN1(n6300), .IN2(n5714), .IN3(n5722), .IN4(n1563), .Q(n1562)
         );
  OA22X1 U1755 ( .IN1(n5702), .IN2(n1564), .IN3(n6146), .IN4(n5701), .Q(n1563)
         );
  AOI22X1 U1756 ( .IN1(\decodedPacket[2][37] ), .IN2(n5693), .IN3(n5688), 
        .IN4(\decodedPacket[1][37] ), .QN(n1564) );
  OA22X1 U1758 ( .IN1(n6320), .IN2(n5747), .IN3(n5753), .IN4(n1566), .Q(n1565)
         );
  OA22X1 U1764 ( .IN1(n6321), .IN2(n5747), .IN3(n5754), .IN4(n1571), .Q(n1570)
         );
  OA22X1 U1770 ( .IN1(n6322), .IN2(n5747), .IN3(n5754), .IN4(n1576), .Q(n1575)
         );
  OA22X1 U1776 ( .IN1(n6323), .IN2(n5747), .IN3(n5754), .IN4(n1581), .Q(n1580)
         );
  OA22X1 U1782 ( .IN1(n6324), .IN2(n5747), .IN3(n5754), .IN4(n1586), .Q(n1585)
         );
  OA22X1 U1788 ( .IN1(n6325), .IN2(n5747), .IN3(n5754), .IN4(n1591), .Q(n1590)
         );
  OA22X1 U1794 ( .IN1(n6326), .IN2(n5747), .IN3(n5755), .IN4(n1596), .Q(n1595)
         );
  OA22X1 U1800 ( .IN1(n6327), .IN2(n5745), .IN3(n5755), .IN4(n1601), .Q(n1600)
         );
  OA22X1 U1806 ( .IN1(n6328), .IN2(n5747), .IN3(n5755), .IN4(n1606), .Q(n1605)
         );
  OA22X1 U1812 ( .IN1(n6329), .IN2(n5747), .IN3(n5755), .IN4(n1611), .Q(n1610)
         );
  OA22X1 U1818 ( .IN1(n6330), .IN2(n5747), .IN3(n5755), .IN4(n1616), .Q(n1615)
         );
  OA22X1 U1824 ( .IN1(n6331), .IN2(n5748), .IN3(n5756), .IN4(n1621), .Q(n1620)
         );
  OA22X1 U1830 ( .IN1(n6332), .IN2(n5748), .IN3(n5756), .IN4(n1626), .Q(n1625)
         );
  OA22X1 U1836 ( .IN1(n6333), .IN2(n5748), .IN3(n5756), .IN4(n1631), .Q(n1630)
         );
  OA22X1 U1842 ( .IN1(n6334), .IN2(n5748), .IN3(n5756), .IN4(n1636), .Q(n1635)
         );
  OA22X1 U1848 ( .IN1(n6335), .IN2(n5748), .IN3(n5756), .IN4(n1641), .Q(n1640)
         );
  OA22X1 U1854 ( .IN1(n6336), .IN2(n5748), .IN3(n5757), .IN4(n1646), .Q(n1645)
         );
  OA22X1 U1860 ( .IN1(n6337), .IN2(n5748), .IN3(n5757), .IN4(n1651), .Q(n1650)
         );
  OA22X1 U1866 ( .IN1(n6338), .IN2(n5748), .IN3(n5757), .IN4(n1656), .Q(n1655)
         );
  OA22X1 U1872 ( .IN1(n6339), .IN2(n5748), .IN3(n5757), .IN4(n1661), .Q(n1660)
         );
  OA22X1 U1878 ( .IN1(n6340), .IN2(n5748), .IN3(n5757), .IN4(n1666), .Q(n1665)
         );
  OA22X1 U1884 ( .IN1(n6341), .IN2(n5748), .IN3(n5753), .IN4(n1671), .Q(n1670)
         );
  OA22X1 U1890 ( .IN1(n6342), .IN2(n5748), .IN3(n5758), .IN4(n1676), .Q(n1675)
         );
  OA22X1 U1896 ( .IN1(n6343), .IN2(n5748), .IN3(n5759), .IN4(n1681), .Q(n1680)
         );
  OA22X1 U1902 ( .IN1(n6344), .IN2(n5748), .IN3(n5755), .IN4(n1686), .Q(n1685)
         );
  OA22X1 U1908 ( .IN1(n6345), .IN2(n5749), .IN3(n5752), .IN4(n1691), .Q(n1690)
         );
  OA22X1 U1914 ( .IN1(n6346), .IN2(n5749), .IN3(n5750), .IN4(n1696), .Q(n1695)
         );
  OA22X1 U1920 ( .IN1(n6315), .IN2(n5749), .IN3(n5751), .IN4(n1701), .Q(n1700)
         );
  OA22X1 U1926 ( .IN1(n6316), .IN2(n5749), .IN3(n5752), .IN4(n1706), .Q(n1705)
         );
  OA22X1 U1932 ( .IN1(n6317), .IN2(n5749), .IN3(n5757), .IN4(n1711), .Q(n1710)
         );
  OA22X1 U1938 ( .IN1(n6318), .IN2(n5749), .IN3(n5756), .IN4(n1716), .Q(n1715)
         );
  OA22X1 U1944 ( .IN1(n6319), .IN2(n5749), .IN3(n5754), .IN4(n1721), .Q(n1720)
         );
  OAI22X1 U1949 ( .IN1(n6455), .IN2(n5772), .IN3(n5765), .IN4(n1725), .QN(
        N9802) );
  OA22X1 U1950 ( .IN1(n6455), .IN2(n5749), .IN3(n5757), .IN4(n1726), .Q(n1725)
         );
  OA22X1 U1951 ( .IN1(n5733), .IN2(n1727), .IN3(n6301), .IN4(n5732), .Q(n1726)
         );
  OA22X1 U1952 ( .IN1(n6301), .IN2(n5716), .IN3(n5722), .IN4(n1728), .Q(n1727)
         );
  OA22X1 U1953 ( .IN1(n5702), .IN2(n1729), .IN3(n6147), .IN4(n5701), .Q(n1728)
         );
  AOI22X1 U1954 ( .IN1(\decodedPacket[2][4] ), .IN2(n5693), .IN3(n5689), .IN4(
        \decodedPacket[1][4] ), .QN(n1729) );
  OAI22X1 U1955 ( .IN1(n6456), .IN2(n5772), .IN3(n5762), .IN4(n1730), .QN(
        N9801) );
  OA22X1 U1956 ( .IN1(n6456), .IN2(n5749), .IN3(n5758), .IN4(n1731), .Q(n1730)
         );
  OA22X1 U1957 ( .IN1(n5733), .IN2(n1732), .IN3(n6302), .IN4(n5732), .Q(n1731)
         );
  OA22X1 U1958 ( .IN1(n6302), .IN2(n5716), .IN3(n5726), .IN4(n1733), .Q(n1732)
         );
  OA22X1 U1959 ( .IN1(n5702), .IN2(n1734), .IN3(n6148), .IN4(n5701), .Q(n1733)
         );
  AOI22X1 U1960 ( .IN1(\decodedPacket[2][3] ), .IN2(n5693), .IN3(n5690), .IN4(
        \decodedPacket[1][3] ), .QN(n1734) );
  OAI22X1 U1961 ( .IN1(n6457), .IN2(n5772), .IN3(n5761), .IN4(n1735), .QN(
        N9800) );
  OA22X1 U1962 ( .IN1(n6457), .IN2(n5749), .IN3(n5751), .IN4(n1736), .Q(n1735)
         );
  OA22X1 U1963 ( .IN1(n5733), .IN2(n1737), .IN3(n6303), .IN4(n5732), .Q(n1736)
         );
  OA22X1 U1964 ( .IN1(n6303), .IN2(n5716), .IN3(n5724), .IN4(n1738), .Q(n1737)
         );
  OA22X1 U1965 ( .IN1(n5702), .IN2(n1739), .IN3(n6149), .IN4(n5701), .Q(n1738)
         );
  AOI22X1 U1966 ( .IN1(\decodedPacket[2][2] ), .IN2(n5693), .IN3(n5683), .IN4(
        \decodedPacket[1][2] ), .QN(n1739) );
  OAI22X1 U1967 ( .IN1(n6458), .IN2(n5772), .IN3(n5762), .IN4(n1740), .QN(
        N9799) );
  OA22X1 U1968 ( .IN1(n6458), .IN2(n5749), .IN3(n5754), .IN4(n1741), .Q(n1740)
         );
  OA22X1 U1969 ( .IN1(n5733), .IN2(n1742), .IN3(n6304), .IN4(n5732), .Q(n1741)
         );
  OA22X1 U1970 ( .IN1(n6304), .IN2(n5716), .IN3(n5725), .IN4(n1743), .Q(n1742)
         );
  OA22X1 U1971 ( .IN1(n5702), .IN2(n1744), .IN3(n6150), .IN4(n5701), .Q(n1743)
         );
  AOI22X1 U1972 ( .IN1(\decodedPacket[2][1] ), .IN2(n5693), .IN3(n5685), .IN4(
        \decodedPacket[1][1] ), .QN(n1744) );
  OAI22X1 U1973 ( .IN1(n6459), .IN2(n5772), .IN3(n5761), .IN4(n1745), .QN(
        N9798) );
  OA22X1 U1974 ( .IN1(n6459), .IN2(n5744), .IN3(n5754), .IN4(n1746), .Q(n1745)
         );
  OA22X1 U1975 ( .IN1(n5733), .IN2(n1747), .IN3(n6305), .IN4(n5732), .Q(n1746)
         );
  OA22X1 U1976 ( .IN1(n6305), .IN2(n5711), .IN3(n5726), .IN4(n1748), .Q(n1747)
         );
  OA22X1 U1977 ( .IN1(n5705), .IN2(n1749), .IN3(n6151), .IN4(n5701), .Q(n1748)
         );
  AOI22X1 U1978 ( .IN1(\decodedPacket[2][0] ), .IN2(n5694), .IN3(n5686), .IN4(
        \decodedPacket[1][0] ), .QN(n1749) );
  NAND4X0 U1979 ( .IN1(n5729), .IN2(n5708), .IN3(n5741), .IN4(n1750), .QN(
        decodedVector_o[1]) );
  NAND4X0 U1981 ( .IN1(n1752), .IN2(decodedPacketValid[7]), .IN3(N8580), .IN4(
        n5987), .QN(n1114) );
  NAND4X0 U1982 ( .IN1(n1753), .IN2(decodedPacketValid[6]), .IN3(N6444), .IN4(
        n5988), .QN(n1116) );
  OA22X1 U2014 ( .IN1(n5653), .IN2(n1788), .IN3(n5856), .IN4(n5666), .Q(n1787)
         );
  OAI22X1 U2020 ( .IN1(n5673), .IN2(n1793), .IN3(n6384), .IN4(n5678), .QN(
        N9791) );
  OA22X1 U2021 ( .IN1(n5653), .IN2(n1794), .IN3(n6349), .IN4(n5663), .Q(n1793)
         );
  OA22X1 U2022 ( .IN1(n6230), .IN2(n5642), .IN3(n5646), .IN4(n1795), .Q(n1794)
         );
  OA22X1 U2023 ( .IN1(n5624), .IN2(n1796), .IN3(n6195), .IN4(n5636), .Q(n1795)
         );
  OA22X1 U2024 ( .IN1(n6076), .IN2(n5621), .IN3(n5622), .IN4(n1797), .Q(n1796)
         );
  OA22X1 U2025 ( .IN1(n5600), .IN2(n1798), .IN3(n6041), .IN4(n5609), .Q(n1797)
         );
  AOI22X1 U2026 ( .IN1(n5591), .IN2(\decodedPacket[1][120] ), .IN3(
        \decodedPacket[0][120] ), .IN4(n5589), .QN(n1798) );
  OAI22X1 U2027 ( .IN1(n5673), .IN2(n1799), .IN3(n6376), .IN4(n5682), .QN(
        N9790) );
  OA22X1 U2028 ( .IN1(n5653), .IN2(n1800), .IN3(n6348), .IN4(n5664), .Q(n1799)
         );
  OA22X1 U2029 ( .IN1(n6222), .IN2(n5642), .IN3(n5647), .IN4(n1801), .Q(n1800)
         );
  OA22X1 U2030 ( .IN1(n5624), .IN2(n1802), .IN3(n6194), .IN4(n5636), .Q(n1801)
         );
  OA22X1 U2031 ( .IN1(n6068), .IN2(n5621), .IN3(n5623), .IN4(n1803), .Q(n1802)
         );
  OA22X1 U2032 ( .IN1(n5600), .IN2(n1804), .IN3(n6040), .IN4(n5610), .Q(n1803)
         );
  AOI22X1 U2033 ( .IN1(n5591), .IN2(\decodedPacket[1][119] ), .IN3(
        \decodedPacket[0][119] ), .IN4(n5588), .QN(n1804) );
  OAI22X1 U2034 ( .IN1(n5673), .IN2(n1805), .IN3(n6373), .IN4(n5680), .QN(
        N9789) );
  OA22X1 U2035 ( .IN1(n5653), .IN2(n1806), .IN3(n6374), .IN4(n5664), .Q(n1805)
         );
  OA22X1 U2036 ( .IN1(n6219), .IN2(n5642), .IN3(n5647), .IN4(n1807), .Q(n1806)
         );
  OA22X1 U2037 ( .IN1(n5624), .IN2(n1808), .IN3(n6220), .IN4(n5636), .Q(n1807)
         );
  OA22X1 U2038 ( .IN1(n6065), .IN2(n5621), .IN3(n5623), .IN4(n1809), .Q(n1808)
         );
  OA22X1 U2039 ( .IN1(n5600), .IN2(n1810), .IN3(n6066), .IN4(n5612), .Q(n1809)
         );
  AOI22X1 U2040 ( .IN1(n5591), .IN2(\decodedPacket[1][118] ), .IN3(
        \decodedPacket[0][118] ), .IN4(n5588), .QN(n1810) );
  OA22X1 U2042 ( .IN1(n5653), .IN2(n1812), .IN3(n6371), .IN4(n5664), .Q(n1811)
         );
  OAI22X1 U2048 ( .IN1(n5673), .IN2(n1817), .IN3(n6373), .IN4(n5681), .QN(
        N9787) );
  OA22X1 U2049 ( .IN1(n5653), .IN2(n1818), .IN3(n6370), .IN4(n5664), .Q(n1817)
         );
  OA22X1 U2050 ( .IN1(n6219), .IN2(n5642), .IN3(n5648), .IN4(n1819), .Q(n1818)
         );
  OA22X1 U2051 ( .IN1(n5624), .IN2(n1820), .IN3(n6216), .IN4(n5636), .Q(n1819)
         );
  OA22X1 U2052 ( .IN1(n6065), .IN2(n5621), .IN3(n5623), .IN4(n1821), .Q(n1820)
         );
  OA22X1 U2053 ( .IN1(n5600), .IN2(n1822), .IN3(n6062), .IN4(n5615), .Q(n1821)
         );
  AOI22X1 U2054 ( .IN1(n5591), .IN2(\decodedPacket[1][116] ), .IN3(
        \decodedPacket[0][116] ), .IN4(n5588), .QN(n1822) );
  OAI22X1 U2055 ( .IN1(n5673), .IN2(n1823), .IN3(n6399), .IN4(n5682), .QN(
        N9786) );
  OA22X1 U2056 ( .IN1(n5653), .IN2(n1824), .IN3(n6347), .IN4(n5664), .Q(n1823)
         );
  OA22X1 U2057 ( .IN1(n6245), .IN2(n5642), .IN3(n5643), .IN4(n1825), .Q(n1824)
         );
  OA22X1 U2058 ( .IN1(n5624), .IN2(n1826), .IN3(n6193), .IN4(n5636), .Q(n1825)
         );
  OA22X1 U2059 ( .IN1(n6091), .IN2(n5621), .IN3(n5623), .IN4(n1827), .Q(n1826)
         );
  OA22X1 U2060 ( .IN1(n5600), .IN2(n1828), .IN3(n6039), .IN4(n5598), .Q(n1827)
         );
  AOI22X1 U2061 ( .IN1(n5591), .IN2(\decodedPacket[1][115] ), .IN3(
        \decodedPacket[0][115] ), .IN4(n5588), .QN(n1828) );
  OAI22X1 U2062 ( .IN1(n5673), .IN2(n1829), .IN3(n5967), .IN4(n5677), .QN(
        N9785) );
  OA22X1 U2063 ( .IN1(n5653), .IN2(n1830), .IN3(n6369), .IN4(n5664), .Q(n1829)
         );
  OA22X1 U2064 ( .IN1(n5952), .IN2(n5642), .IN3(n5643), .IN4(n1831), .Q(n1830)
         );
  OA22X1 U2065 ( .IN1(n5624), .IN2(n1832), .IN3(n6215), .IN4(n5636), .Q(n1831)
         );
  OA22X1 U2066 ( .IN1(n5937), .IN2(n5621), .IN3(n5623), .IN4(n1833), .Q(n1832)
         );
  OA22X1 U2067 ( .IN1(n5600), .IN2(n1834), .IN3(n6061), .IN4(n5598), .Q(n1833)
         );
  AOI22X1 U2068 ( .IN1(n5591), .IN2(\decodedPacket[1][114] ), .IN3(
        \decodedPacket[0][114] ), .IN4(n5588), .QN(n1834) );
  OAI22X1 U2069 ( .IN1(n5674), .IN2(n1835), .IN3(n5968), .IN4(n5680), .QN(
        N9784) );
  OA22X1 U2070 ( .IN1(n5653), .IN2(n1836), .IN3(n6368), .IN4(n5664), .Q(n1835)
         );
  OA22X1 U2071 ( .IN1(n5953), .IN2(n5642), .IN3(n5643), .IN4(n1837), .Q(n1836)
         );
  OA22X1 U2072 ( .IN1(n5624), .IN2(n1838), .IN3(n6214), .IN4(n5636), .Q(n1837)
         );
  OA22X1 U2073 ( .IN1(n5938), .IN2(n5621), .IN3(n5623), .IN4(n1839), .Q(n1838)
         );
  OA22X1 U2074 ( .IN1(n5600), .IN2(n1840), .IN3(n6060), .IN4(n5597), .Q(n1839)
         );
  AOI22X1 U2075 ( .IN1(n5591), .IN2(\decodedPacket[1][113] ), .IN3(
        \decodedPacket[0][113] ), .IN4(n5588), .QN(n1840) );
  OAI22X1 U2076 ( .IN1(n5674), .IN2(n1841), .IN3(n5969), .IN4(n5682), .QN(
        N9783) );
  OA22X1 U2077 ( .IN1(n5653), .IN2(n1842), .IN3(n6367), .IN4(n5664), .Q(n1841)
         );
  OA22X1 U2078 ( .IN1(n5954), .IN2(n5642), .IN3(n5643), .IN4(n1843), .Q(n1842)
         );
  OA22X1 U2079 ( .IN1(n5624), .IN2(n1844), .IN3(n6213), .IN4(n5635), .Q(n1843)
         );
  OA22X1 U2080 ( .IN1(n5939), .IN2(n5621), .IN3(n5623), .IN4(n1845), .Q(n1844)
         );
  OA22X1 U2081 ( .IN1(n5600), .IN2(n1846), .IN3(n6059), .IN4(n5614), .Q(n1845)
         );
  AOI22X1 U2082 ( .IN1(n5591), .IN2(\decodedPacket[1][112] ), .IN3(
        \decodedPacket[0][112] ), .IN4(n5588), .QN(n1846) );
  OAI22X1 U2083 ( .IN1(n5674), .IN2(n1847), .IN3(n5970), .IN4(n5680), .QN(
        N9782) );
  OA22X1 U2084 ( .IN1(n5653), .IN2(n1848), .IN3(n6366), .IN4(n5664), .Q(n1847)
         );
  OA22X1 U2085 ( .IN1(n5955), .IN2(n5642), .IN3(n5643), .IN4(n1849), .Q(n1848)
         );
  OA22X1 U2086 ( .IN1(n5624), .IN2(n1850), .IN3(n6212), .IN4(n5635), .Q(n1849)
         );
  OA22X1 U2087 ( .IN1(n5940), .IN2(n5621), .IN3(n5623), .IN4(n1851), .Q(n1850)
         );
  OA22X1 U2088 ( .IN1(n5600), .IN2(n1852), .IN3(n6058), .IN4(n5615), .Q(n1851)
         );
  AOI22X1 U2089 ( .IN1(n5591), .IN2(\decodedPacket[1][111] ), .IN3(
        \decodedPacket[0][111] ), .IN4(n5589), .QN(n1852) );
  OAI22X1 U2090 ( .IN1(n5674), .IN2(n1853), .IN3(n5971), .IN4(n5680), .QN(
        N9781) );
  OA22X1 U2091 ( .IN1(n5653), .IN2(n1854), .IN3(n6365), .IN4(n5664), .Q(n1853)
         );
  OA22X1 U2092 ( .IN1(n5956), .IN2(n5642), .IN3(n5644), .IN4(n1855), .Q(n1854)
         );
  OA22X1 U2093 ( .IN1(n5624), .IN2(n1856), .IN3(n6211), .IN4(n5635), .Q(n1855)
         );
  OA22X1 U2094 ( .IN1(n5941), .IN2(n5621), .IN3(n5623), .IN4(n1857), .Q(n1856)
         );
  OA22X1 U2095 ( .IN1(n5600), .IN2(n1858), .IN3(n6057), .IN4(n5615), .Q(n1857)
         );
  AOI22X1 U2096 ( .IN1(n5591), .IN2(\decodedPacket[1][110] ), .IN3(
        \decodedPacket[0][110] ), .IN4(n5589), .QN(n1858) );
  OAI22X1 U2097 ( .IN1(n5674), .IN2(n1859), .IN3(n5972), .IN4(n5682), .QN(
        N9780) );
  OA22X1 U2098 ( .IN1(n5654), .IN2(n1860), .IN3(n6364), .IN4(n5664), .Q(n1859)
         );
  OA22X1 U2099 ( .IN1(n5957), .IN2(n5642), .IN3(n5644), .IN4(n1861), .Q(n1860)
         );
  OA22X1 U2100 ( .IN1(n5624), .IN2(n1862), .IN3(n6210), .IN4(n5635), .Q(n1861)
         );
  OA22X1 U2101 ( .IN1(n5942), .IN2(n5621), .IN3(n5623), .IN4(n1863), .Q(n1862)
         );
  OA22X1 U2102 ( .IN1(n5600), .IN2(n1864), .IN3(n6056), .IN4(n5615), .Q(n1863)
         );
  AOI22X1 U2103 ( .IN1(n5592), .IN2(\decodedPacket[1][109] ), .IN3(
        \decodedPacket[0][109] ), .IN4(n5589), .QN(n1864) );
  OAI22X1 U2104 ( .IN1(n5674), .IN2(n1865), .IN3(n5973), .IN4(n5681), .QN(
        N9779) );
  OA22X1 U2105 ( .IN1(n5654), .IN2(n1866), .IN3(n6363), .IN4(n5664), .Q(n1865)
         );
  OA22X1 U2106 ( .IN1(n5958), .IN2(n5642), .IN3(n5644), .IN4(n1867), .Q(n1866)
         );
  OA22X1 U2107 ( .IN1(n5624), .IN2(n1868), .IN3(n6209), .IN4(n5635), .Q(n1867)
         );
  OA22X1 U2108 ( .IN1(n5943), .IN2(n5621), .IN3(n5623), .IN4(n1869), .Q(n1868)
         );
  OA22X1 U2109 ( .IN1(n5600), .IN2(n1870), .IN3(n6055), .IN4(n5615), .Q(n1869)
         );
  AOI22X1 U2110 ( .IN1(n5592), .IN2(\decodedPacket[1][108] ), .IN3(
        \decodedPacket[0][108] ), .IN4(n5589), .QN(n1870) );
  OAI22X1 U2111 ( .IN1(n5674), .IN2(n1871), .IN3(n5974), .IN4(n5676), .QN(
        N9778) );
  OA22X1 U2112 ( .IN1(n5654), .IN2(n1872), .IN3(n6362), .IN4(n5664), .Q(n1871)
         );
  OA22X1 U2113 ( .IN1(n5959), .IN2(n5642), .IN3(n5644), .IN4(n1873), .Q(n1872)
         );
  OA22X1 U2114 ( .IN1(n5624), .IN2(n1874), .IN3(n6208), .IN4(n5635), .Q(n1873)
         );
  OA22X1 U2115 ( .IN1(n5944), .IN2(n5621), .IN3(n5623), .IN4(n1875), .Q(n1874)
         );
  OA22X1 U2116 ( .IN1(n5601), .IN2(n1876), .IN3(n6054), .IN4(n5615), .Q(n1875)
         );
  AOI22X1 U2117 ( .IN1(n5592), .IN2(\decodedPacket[1][107] ), .IN3(
        \decodedPacket[0][107] ), .IN4(n5589), .QN(n1876) );
  OAI22X1 U2118 ( .IN1(n5674), .IN2(n1877), .IN3(n5975), .IN4(n1757), .QN(
        N9777) );
  OA22X1 U2119 ( .IN1(n5654), .IN2(n1878), .IN3(n6308), .IN4(n5664), .Q(n1877)
         );
  OA22X1 U2120 ( .IN1(n5960), .IN2(n5642), .IN3(n5644), .IN4(n1879), .Q(n1878)
         );
  OA22X1 U2121 ( .IN1(n5624), .IN2(n1880), .IN3(n6154), .IN4(n5635), .Q(n1879)
         );
  OA22X1 U2122 ( .IN1(n5945), .IN2(n5621), .IN3(n5623), .IN4(n1881), .Q(n1880)
         );
  OA22X1 U2123 ( .IN1(n5601), .IN2(n1882), .IN3(n6000), .IN4(n5615), .Q(n1881)
         );
  AOI22X1 U2124 ( .IN1(n5592), .IN2(\decodedPacket[1][106] ), .IN3(
        \decodedPacket[0][106] ), .IN4(n5589), .QN(n1882) );
  OAI22X1 U2125 ( .IN1(n5674), .IN2(n1883), .IN3(n5976), .IN4(n5681), .QN(
        N9776) );
  OA22X1 U2126 ( .IN1(n5654), .IN2(n1884), .IN3(n6309), .IN4(n5664), .Q(n1883)
         );
  OA22X1 U2127 ( .IN1(n5961), .IN2(n5642), .IN3(n5645), .IN4(n1885), .Q(n1884)
         );
  OA22X1 U2128 ( .IN1(n5624), .IN2(n1886), .IN3(n6155), .IN4(n5635), .Q(n1885)
         );
  OA22X1 U2129 ( .IN1(n5946), .IN2(n5621), .IN3(n5623), .IN4(n1887), .Q(n1886)
         );
  OA22X1 U2130 ( .IN1(n5601), .IN2(n1888), .IN3(n6001), .IN4(n5614), .Q(n1887)
         );
  AOI22X1 U2131 ( .IN1(n5592), .IN2(\decodedPacket[1][105] ), .IN3(
        \decodedPacket[0][105] ), .IN4(n5589), .QN(n1888) );
  OAI22X1 U2132 ( .IN1(n5674), .IN2(n1889), .IN3(n5977), .IN4(n5679), .QN(
        N9775) );
  OA22X1 U2133 ( .IN1(n5654), .IN2(n1890), .IN3(n6310), .IN4(n5652), .Q(n1889)
         );
  OA22X1 U2134 ( .IN1(n5962), .IN2(n5642), .IN3(n5645), .IN4(n1891), .Q(n1890)
         );
  OA22X1 U2135 ( .IN1(n5624), .IN2(n1892), .IN3(n6156), .IN4(n5635), .Q(n1891)
         );
  OA22X1 U2136 ( .IN1(n5947), .IN2(n5621), .IN3(n5623), .IN4(n1893), .Q(n1892)
         );
  OA22X1 U2137 ( .IN1(n5601), .IN2(n1894), .IN3(n6002), .IN4(n5614), .Q(n1893)
         );
  AOI22X1 U2138 ( .IN1(n5592), .IN2(\decodedPacket[1][104] ), .IN3(
        \decodedPacket[0][104] ), .IN4(n5589), .QN(n1894) );
  OAI22X1 U2139 ( .IN1(n5674), .IN2(n1895), .IN3(n5978), .IN4(n5677), .QN(
        N9774) );
  OA22X1 U2140 ( .IN1(n5654), .IN2(n1896), .IN3(n6311), .IN4(n5651), .Q(n1895)
         );
  OA22X1 U2141 ( .IN1(n5963), .IN2(n5642), .IN3(n5645), .IN4(n1897), .Q(n1896)
         );
  OA22X1 U2142 ( .IN1(n5624), .IN2(n1898), .IN3(n6157), .IN4(n5635), .Q(n1897)
         );
  OA22X1 U2143 ( .IN1(n5948), .IN2(n5620), .IN3(n5623), .IN4(n1899), .Q(n1898)
         );
  OA22X1 U2144 ( .IN1(n5601), .IN2(n1900), .IN3(n6003), .IN4(n5614), .Q(n1899)
         );
  AOI22X1 U2145 ( .IN1(n5592), .IN2(\decodedPacket[1][103] ), .IN3(
        \decodedPacket[0][103] ), .IN4(n5589), .QN(n1900) );
  OAI22X1 U2146 ( .IN1(n5674), .IN2(n1901), .IN3(n5979), .IN4(n5679), .QN(
        N9773) );
  OA22X1 U2147 ( .IN1(n5654), .IN2(n1902), .IN3(n6312), .IN4(n5652), .Q(n1901)
         );
  OA22X1 U2148 ( .IN1(n5964), .IN2(n5641), .IN3(n5645), .IN4(n1903), .Q(n1902)
         );
  OA22X1 U2149 ( .IN1(n5624), .IN2(n1904), .IN3(n6158), .IN4(n5635), .Q(n1903)
         );
  OA22X1 U2150 ( .IN1(n5949), .IN2(n5620), .IN3(n5623), .IN4(n1905), .Q(n1904)
         );
  OA22X1 U2151 ( .IN1(n5601), .IN2(n1906), .IN3(n6004), .IN4(n5614), .Q(n1905)
         );
  AOI22X1 U2152 ( .IN1(n5592), .IN2(\decodedPacket[1][102] ), .IN3(
        \decodedPacket[0][102] ), .IN4(n5589), .QN(n1906) );
  OAI22X1 U2153 ( .IN1(n5674), .IN2(n1907), .IN3(n5980), .IN4(n5682), .QN(
        N9772) );
  OA22X1 U2154 ( .IN1(n5654), .IN2(n1908), .IN3(n6313), .IN4(n5651), .Q(n1907)
         );
  OA22X1 U2155 ( .IN1(n5965), .IN2(n5641), .IN3(n5645), .IN4(n1909), .Q(n1908)
         );
  OA22X1 U2156 ( .IN1(n5624), .IN2(n1910), .IN3(n6159), .IN4(n5635), .Q(n1909)
         );
  OA22X1 U2157 ( .IN1(n5950), .IN2(n5620), .IN3(n5623), .IN4(n1911), .Q(n1910)
         );
  OA22X1 U2158 ( .IN1(n5601), .IN2(n1912), .IN3(n6005), .IN4(n5614), .Q(n1911)
         );
  AOI22X1 U2159 ( .IN1(n5592), .IN2(\decodedPacket[1][101] ), .IN3(
        \decodedPacket[0][101] ), .IN4(n5589), .QN(n1912) );
  OAI22X1 U2160 ( .IN1(n5674), .IN2(n1913), .IN3(n5981), .IN4(n5678), .QN(
        N9771) );
  OA22X1 U2161 ( .IN1(n5654), .IN2(n1914), .IN3(n6314), .IN4(n5652), .Q(n1913)
         );
  OA22X1 U2162 ( .IN1(n5966), .IN2(n5641), .IN3(n5646), .IN4(n1915), .Q(n1914)
         );
  OA22X1 U2163 ( .IN1(n5624), .IN2(n1916), .IN3(n6160), .IN4(n5635), .Q(n1915)
         );
  OA22X1 U2164 ( .IN1(n5951), .IN2(n5620), .IN3(n5623), .IN4(n1917), .Q(n1916)
         );
  OA22X1 U2165 ( .IN1(n5601), .IN2(n1918), .IN3(n6006), .IN4(n5613), .Q(n1917)
         );
  AOI22X1 U2166 ( .IN1(n5592), .IN2(\decodedPacket[1][100] ), .IN3(
        \decodedPacket[0][100] ), .IN4(n5589), .QN(n1918) );
  OAI22X1 U2167 ( .IN1(n5674), .IN2(n1919), .IN3(n6375), .IN4(n5679), .QN(
        N9770) );
  OA22X1 U2168 ( .IN1(n5654), .IN2(n1920), .IN3(n6307), .IN4(n5651), .Q(n1919)
         );
  OA22X1 U2169 ( .IN1(n6221), .IN2(n5641), .IN3(n5649), .IN4(n1921), .Q(n1920)
         );
  OA22X1 U2170 ( .IN1(n5624), .IN2(n1922), .IN3(n6153), .IN4(n5634), .Q(n1921)
         );
  OA22X1 U2171 ( .IN1(n6067), .IN2(n5620), .IN3(n5623), .IN4(n1923), .Q(n1922)
         );
  OA22X1 U2172 ( .IN1(n5601), .IN2(n1924), .IN3(n5999), .IN4(n5613), .Q(n1923)
         );
  AOI22X1 U2173 ( .IN1(n5592), .IN2(\decodedPacket[1][99] ), .IN3(
        \decodedPacket[0][99] ), .IN4(n5589), .QN(n1924) );
  OAI22X1 U2174 ( .IN1(n5674), .IN2(n1925), .IN3(n6372), .IN4(n1757), .QN(
        N9769) );
  OA22X1 U2175 ( .IN1(n5654), .IN2(n1926), .IN3(n6306), .IN4(n5652), .Q(n1925)
         );
  OA22X1 U2176 ( .IN1(n6218), .IN2(n5641), .IN3(n5645), .IN4(n1927), .Q(n1926)
         );
  OA22X1 U2177 ( .IN1(n5624), .IN2(n1928), .IN3(n6152), .IN4(n5634), .Q(n1927)
         );
  OA22X1 U2178 ( .IN1(n6064), .IN2(n5620), .IN3(n5623), .IN4(n1929), .Q(n1928)
         );
  OA22X1 U2179 ( .IN1(n5601), .IN2(n1930), .IN3(n5998), .IN4(n5613), .Q(n1929)
         );
  AOI22X1 U2180 ( .IN1(n5592), .IN2(\decodedPacket[1][98] ), .IN3(
        \decodedPacket[0][98] ), .IN4(n5589), .QN(n1930) );
  OAI22X1 U2181 ( .IN1(n5674), .IN2(n1931), .IN3(n6377), .IN4(n5681), .QN(
        N9768) );
  OA22X1 U2182 ( .IN1(n5655), .IN2(n1932), .IN3(n6422), .IN4(n5651), .Q(n1931)
         );
  OA22X1 U2183 ( .IN1(n6223), .IN2(n5641), .IN3(n5648), .IN4(n1933), .Q(n1932)
         );
  OA22X1 U2184 ( .IN1(n5624), .IN2(n1934), .IN3(n6268), .IN4(n5634), .Q(n1933)
         );
  OA22X1 U2185 ( .IN1(n6069), .IN2(n5620), .IN3(n5623), .IN4(n1935), .Q(n1934)
         );
  OA22X1 U2186 ( .IN1(n5601), .IN2(n1936), .IN3(n6114), .IN4(n5613), .Q(n1935)
         );
  AOI22X1 U2187 ( .IN1(n5592), .IN2(\decodedPacket[1][97] ), .IN3(
        \decodedPacket[0][97] ), .IN4(n5589), .QN(n1936) );
  OAI22X1 U2188 ( .IN1(n5674), .IN2(n1937), .IN3(n6378), .IN4(n5682), .QN(
        N9766) );
  OA22X1 U2189 ( .IN1(n5655), .IN2(n1938), .IN3(n6421), .IN4(n5652), .Q(n1937)
         );
  OA22X1 U2190 ( .IN1(n6224), .IN2(n5641), .IN3(n5650), .IN4(n1939), .Q(n1938)
         );
  OA22X1 U2191 ( .IN1(n5624), .IN2(n1940), .IN3(n6267), .IN4(n5634), .Q(n1939)
         );
  OA22X1 U2192 ( .IN1(n6070), .IN2(n5620), .IN3(n5623), .IN4(n1941), .Q(n1940)
         );
  OA22X1 U2193 ( .IN1(n5601), .IN2(n1942), .IN3(n6113), .IN4(n5613), .Q(n1941)
         );
  AOI22X1 U2194 ( .IN1(n5592), .IN2(\decodedPacket[1][96] ), .IN3(
        \decodedPacket[0][96] ), .IN4(n5589), .QN(n1942) );
  OAI22X1 U2195 ( .IN1(n5674), .IN2(n1943), .IN3(n6379), .IN4(n5682), .QN(
        N9765) );
  OA22X1 U2196 ( .IN1(n5655), .IN2(n1944), .IN3(n6420), .IN4(n5651), .Q(n1943)
         );
  OA22X1 U2197 ( .IN1(n6225), .IN2(n5641), .IN3(n5650), .IN4(n1945), .Q(n1944)
         );
  OA22X1 U2198 ( .IN1(n5624), .IN2(n1946), .IN3(n6266), .IN4(n5634), .Q(n1945)
         );
  OA22X1 U2199 ( .IN1(n6071), .IN2(n5620), .IN3(n5623), .IN4(n1947), .Q(n1946)
         );
  OA22X1 U2200 ( .IN1(n5601), .IN2(n1948), .IN3(n6112), .IN4(n5609), .Q(n1947)
         );
  AOI22X1 U2201 ( .IN1(n5592), .IN2(\decodedPacket[1][95] ), .IN3(
        \decodedPacket[0][95] ), .IN4(n5589), .QN(n1948) );
  OAI22X1 U2202 ( .IN1(n5674), .IN2(n1949), .IN3(n6380), .IN4(n5682), .QN(
        N9764) );
  OA22X1 U2203 ( .IN1(n5655), .IN2(n1950), .IN3(n6419), .IN4(n5652), .Q(n1949)
         );
  OA22X1 U2204 ( .IN1(n6226), .IN2(n5641), .IN3(n5647), .IN4(n1951), .Q(n1950)
         );
  OA22X1 U2205 ( .IN1(n5624), .IN2(n1952), .IN3(n6265), .IN4(n5634), .Q(n1951)
         );
  OA22X1 U2206 ( .IN1(n6072), .IN2(n5620), .IN3(n5623), .IN4(n1953), .Q(n1952)
         );
  OA22X1 U2207 ( .IN1(n5601), .IN2(n1954), .IN3(n6111), .IN4(n5610), .Q(n1953)
         );
  AOI22X1 U2208 ( .IN1(n5592), .IN2(\decodedPacket[1][94] ), .IN3(
        \decodedPacket[0][94] ), .IN4(n5589), .QN(n1954) );
  OAI22X1 U2209 ( .IN1(n5674), .IN2(n1955), .IN3(n6381), .IN4(n5682), .QN(
        N9763) );
  OA22X1 U2210 ( .IN1(n5655), .IN2(n1956), .IN3(n6418), .IN4(n5651), .Q(n1955)
         );
  OA22X1 U2211 ( .IN1(n6227), .IN2(n5641), .IN3(n5643), .IN4(n1957), .Q(n1956)
         );
  OA22X1 U2212 ( .IN1(n5624), .IN2(n1958), .IN3(n6264), .IN4(n5634), .Q(n1957)
         );
  OA22X1 U2213 ( .IN1(n6073), .IN2(n5620), .IN3(n5623), .IN4(n1959), .Q(n1958)
         );
  OA22X1 U2214 ( .IN1(n5601), .IN2(n1960), .IN3(n6110), .IN4(n5612), .Q(n1959)
         );
  AOI22X1 U2215 ( .IN1(n5592), .IN2(\decodedPacket[1][93] ), .IN3(
        \decodedPacket[0][93] ), .IN4(n5589), .QN(n1960) );
  OAI22X1 U2216 ( .IN1(n5674), .IN2(n1961), .IN3(n6382), .IN4(n5682), .QN(
        N9762) );
  OA22X1 U2217 ( .IN1(n5655), .IN2(n1962), .IN3(n6417), .IN4(n5652), .Q(n1961)
         );
  OA22X1 U2218 ( .IN1(n6228), .IN2(n5641), .IN3(n5644), .IN4(n1963), .Q(n1962)
         );
  OA22X1 U2219 ( .IN1(n5624), .IN2(n1964), .IN3(n6263), .IN4(n5634), .Q(n1963)
         );
  OA22X1 U2220 ( .IN1(n6074), .IN2(n5620), .IN3(n5623), .IN4(n1965), .Q(n1964)
         );
  OA22X1 U2221 ( .IN1(n5602), .IN2(n1966), .IN3(n6109), .IN4(n5612), .Q(n1965)
         );
  AOI22X1 U2222 ( .IN1(n5593), .IN2(\decodedPacket[1][92] ), .IN3(
        \decodedPacket[0][92] ), .IN4(n5589), .QN(n1966) );
  OAI22X1 U2223 ( .IN1(n5674), .IN2(n1967), .IN3(n6383), .IN4(n5682), .QN(
        N9761) );
  OA22X1 U2224 ( .IN1(n5655), .IN2(n1968), .IN3(n6416), .IN4(n5651), .Q(n1967)
         );
  OA22X1 U2225 ( .IN1(n6229), .IN2(n5641), .IN3(n5646), .IN4(n1969), .Q(n1968)
         );
  OA22X1 U2226 ( .IN1(n5624), .IN2(n1970), .IN3(n6262), .IN4(n5634), .Q(n1969)
         );
  OA22X1 U2227 ( .IN1(n6075), .IN2(n5620), .IN3(n5623), .IN4(n1971), .Q(n1970)
         );
  OA22X1 U2228 ( .IN1(n5602), .IN2(n1972), .IN3(n6108), .IN4(n5599), .Q(n1971)
         );
  AOI22X1 U2229 ( .IN1(n5593), .IN2(\decodedPacket[1][91] ), .IN3(
        \decodedPacket[0][91] ), .IN4(n5589), .QN(n1972) );
  OAI22X1 U2230 ( .IN1(n5674), .IN2(n1973), .IN3(n6385), .IN4(n5681), .QN(
        N9760) );
  OA22X1 U2231 ( .IN1(n5655), .IN2(n1974), .IN3(n6359), .IN4(n5652), .Q(n1973)
         );
  OA22X1 U2232 ( .IN1(n6231), .IN2(n5641), .IN3(n5650), .IN4(n1975), .Q(n1974)
         );
  OA22X1 U2233 ( .IN1(n5625), .IN2(n1976), .IN3(n6205), .IN4(n5634), .Q(n1975)
         );
  OA22X1 U2234 ( .IN1(n6077), .IN2(n5620), .IN3(n5623), .IN4(n1977), .Q(n1976)
         );
  OA22X1 U2235 ( .IN1(n5602), .IN2(n1978), .IN3(n6051), .IN4(n5608), .Q(n1977)
         );
  AOI22X1 U2236 ( .IN1(n5593), .IN2(\decodedPacket[1][90] ), .IN3(
        \decodedPacket[0][90] ), .IN4(n5589), .QN(n1978) );
  OAI22X1 U2237 ( .IN1(n5674), .IN2(n1979), .IN3(n6386), .IN4(n5681), .QN(
        N9759) );
  OA22X1 U2238 ( .IN1(n5655), .IN2(n1980), .IN3(n6358), .IN4(n5665), .Q(n1979)
         );
  OA22X1 U2239 ( .IN1(n6232), .IN2(n5641), .IN3(n5647), .IN4(n1981), .Q(n1980)
         );
  OA22X1 U2240 ( .IN1(n5625), .IN2(n1982), .IN3(n6204), .IN4(n5634), .Q(n1981)
         );
  OA22X1 U2241 ( .IN1(n6078), .IN2(n5620), .IN3(n5623), .IN4(n1983), .Q(n1982)
         );
  OA22X1 U2242 ( .IN1(n5602), .IN2(n1984), .IN3(n6050), .IN4(n5611), .Q(n1983)
         );
  AOI22X1 U2243 ( .IN1(n5593), .IN2(\decodedPacket[1][89] ), .IN3(
        \decodedPacket[0][89] ), .IN4(n5589), .QN(n1984) );
  OAI22X1 U2244 ( .IN1(n5674), .IN2(n1985), .IN3(n6387), .IN4(n5681), .QN(
        N9758) );
  OA22X1 U2245 ( .IN1(n5655), .IN2(n1986), .IN3(n6357), .IN4(n5665), .Q(n1985)
         );
  OA22X1 U2246 ( .IN1(n6233), .IN2(n5641), .IN3(n5646), .IN4(n1987), .Q(n1986)
         );
  OA22X1 U2247 ( .IN1(n5625), .IN2(n1988), .IN3(n6203), .IN4(n5634), .Q(n1987)
         );
  OA22X1 U2248 ( .IN1(n6079), .IN2(n5620), .IN3(n5623), .IN4(n1989), .Q(n1988)
         );
  OA22X1 U2249 ( .IN1(n5602), .IN2(n1990), .IN3(n6049), .IN4(n5598), .Q(n1989)
         );
  AOI22X1 U2250 ( .IN1(n5593), .IN2(\decodedPacket[1][88] ), .IN3(
        \decodedPacket[0][88] ), .IN4(n5589), .QN(n1990) );
  OAI22X1 U2251 ( .IN1(n5674), .IN2(n1991), .IN3(n6388), .IN4(n5681), .QN(
        N9757) );
  OA22X1 U2252 ( .IN1(n5655), .IN2(n1992), .IN3(n6356), .IN4(n5665), .Q(n1991)
         );
  OA22X1 U2253 ( .IN1(n6234), .IN2(n5641), .IN3(n5644), .IN4(n1993), .Q(n1992)
         );
  OA22X1 U2254 ( .IN1(n5625), .IN2(n1994), .IN3(n6202), .IN4(n5634), .Q(n1993)
         );
  OA22X1 U2255 ( .IN1(n6080), .IN2(n5620), .IN3(n5623), .IN4(n1995), .Q(n1994)
         );
  OA22X1 U2256 ( .IN1(n5602), .IN2(n1996), .IN3(n6048), .IN4(n5609), .Q(n1995)
         );
  AOI22X1 U2257 ( .IN1(n5593), .IN2(\decodedPacket[1][87] ), .IN3(
        \decodedPacket[0][87] ), .IN4(n5589), .QN(n1996) );
  OAI22X1 U2258 ( .IN1(n5674), .IN2(n1997), .IN3(n6389), .IN4(n5681), .QN(
        N9756) );
  OA22X1 U2259 ( .IN1(n5655), .IN2(n1998), .IN3(n6355), .IN4(n5665), .Q(n1997)
         );
  OA22X1 U2260 ( .IN1(n6235), .IN2(n5641), .IN3(n5649), .IN4(n1999), .Q(n1998)
         );
  OA22X1 U2261 ( .IN1(n5625), .IN2(n2000), .IN3(n6201), .IN4(n5633), .Q(n1999)
         );
  OA22X1 U2262 ( .IN1(n6081), .IN2(n5620), .IN3(n5623), .IN4(n2001), .Q(n2000)
         );
  OA22X1 U2263 ( .IN1(n5602), .IN2(n2002), .IN3(n6047), .IN4(n5610), .Q(n2001)
         );
  AOI22X1 U2264 ( .IN1(n5593), .IN2(\decodedPacket[1][86] ), .IN3(
        \decodedPacket[0][86] ), .IN4(n5589), .QN(n2002) );
  OAI22X1 U2265 ( .IN1(n5674), .IN2(n2003), .IN3(n6390), .IN4(n5681), .QN(
        N9755) );
  OA22X1 U2266 ( .IN1(n5656), .IN2(n2004), .IN3(n6354), .IN4(n5665), .Q(n2003)
         );
  OA22X1 U2267 ( .IN1(n6236), .IN2(n5641), .IN3(n5643), .IN4(n2005), .Q(n2004)
         );
  OA22X1 U2268 ( .IN1(n5625), .IN2(n2006), .IN3(n6200), .IN4(n5633), .Q(n2005)
         );
  OA22X1 U2269 ( .IN1(n6082), .IN2(n5620), .IN3(n5623), .IN4(n2007), .Q(n2006)
         );
  OA22X1 U2270 ( .IN1(n5602), .IN2(n2008), .IN3(n6046), .IN4(n5612), .Q(n2007)
         );
  AOI22X1 U2271 ( .IN1(n5593), .IN2(\decodedPacket[1][85] ), .IN3(
        \decodedPacket[0][85] ), .IN4(n5589), .QN(n2008) );
  OAI22X1 U2272 ( .IN1(n5674), .IN2(n2009), .IN3(n6391), .IN4(n5680), .QN(
        N9754) );
  OA22X1 U2273 ( .IN1(n5656), .IN2(n2010), .IN3(n6353), .IN4(n5665), .Q(n2009)
         );
  OA22X1 U2274 ( .IN1(n6237), .IN2(n5641), .IN3(n5646), .IN4(n2011), .Q(n2010)
         );
  OA22X1 U2275 ( .IN1(n5625), .IN2(n2012), .IN3(n6199), .IN4(n5633), .Q(n2011)
         );
  OA22X1 U2276 ( .IN1(n6083), .IN2(n5620), .IN3(n5623), .IN4(n2013), .Q(n2012)
         );
  OA22X1 U2277 ( .IN1(n5602), .IN2(n2014), .IN3(n6045), .IN4(n5612), .Q(n2013)
         );
  AOI22X1 U2278 ( .IN1(n5593), .IN2(\decodedPacket[1][84] ), .IN3(
        \decodedPacket[0][84] ), .IN4(n5589), .QN(n2014) );
  OAI22X1 U2279 ( .IN1(n5674), .IN2(n2015), .IN3(n6400), .IN4(n5680), .QN(
        N9753) );
  OA22X1 U2280 ( .IN1(n5656), .IN2(n2016), .IN3(n6415), .IN4(n5665), .Q(n2015)
         );
  OA22X1 U2281 ( .IN1(n6246), .IN2(n5641), .IN3(n5644), .IN4(n2017), .Q(n2016)
         );
  OA22X1 U2282 ( .IN1(n5625), .IN2(n2018), .IN3(n6261), .IN4(n5633), .Q(n2017)
         );
  OA22X1 U2283 ( .IN1(n6092), .IN2(n5620), .IN3(n5623), .IN4(n2019), .Q(n2018)
         );
  OA22X1 U2284 ( .IN1(n5602), .IN2(n2020), .IN3(n6107), .IN4(n5612), .Q(n2019)
         );
  AOI22X1 U2285 ( .IN1(n5593), .IN2(\decodedPacket[1][83] ), .IN3(
        \decodedPacket[0][83] ), .IN4(n5589), .QN(n2020) );
  OAI22X1 U2286 ( .IN1(n5674), .IN2(n2021), .IN3(n6406), .IN4(n5680), .QN(
        N9752) );
  OA22X1 U2287 ( .IN1(n5656), .IN2(n2022), .IN3(n6414), .IN4(n5665), .Q(n2021)
         );
  OA22X1 U2288 ( .IN1(n6252), .IN2(n5641), .IN3(n5649), .IN4(n2023), .Q(n2022)
         );
  OA22X1 U2289 ( .IN1(n5625), .IN2(n2024), .IN3(n6260), .IN4(n5633), .Q(n2023)
         );
  OA22X1 U2290 ( .IN1(n6098), .IN2(n5620), .IN3(n5623), .IN4(n2025), .Q(n2024)
         );
  OA22X1 U2291 ( .IN1(n5602), .IN2(n2026), .IN3(n6106), .IN4(n5612), .Q(n2025)
         );
  AOI22X1 U2292 ( .IN1(n5593), .IN2(\decodedPacket[1][82] ), .IN3(
        \decodedPacket[0][82] ), .IN4(n5589), .QN(n2026) );
  OAI22X1 U2293 ( .IN1(n5674), .IN2(n2027), .IN3(n6407), .IN4(n5680), .QN(
        N9751) );
  OA22X1 U2294 ( .IN1(n5656), .IN2(n2028), .IN3(n6413), .IN4(n5665), .Q(n2027)
         );
  OA22X1 U2295 ( .IN1(n6253), .IN2(n5641), .IN3(n5643), .IN4(n2029), .Q(n2028)
         );
  OA22X1 U2296 ( .IN1(n5625), .IN2(n2030), .IN3(n6259), .IN4(n5633), .Q(n2029)
         );
  OA22X1 U2297 ( .IN1(n6099), .IN2(n5620), .IN3(n5623), .IN4(n2031), .Q(n2030)
         );
  OA22X1 U2298 ( .IN1(n5602), .IN2(n2032), .IN3(n6105), .IN4(n5612), .Q(n2031)
         );
  AOI22X1 U2299 ( .IN1(n5593), .IN2(\decodedPacket[1][81] ), .IN3(
        \decodedPacket[0][81] ), .IN4(n5589), .QN(n2032) );
  OAI22X1 U2300 ( .IN1(n5674), .IN2(n2033), .IN3(n6408), .IN4(n5680), .QN(
        N9750) );
  OA22X1 U2301 ( .IN1(n5656), .IN2(n2034), .IN3(n6412), .IN4(n5665), .Q(n2033)
         );
  OA22X1 U2302 ( .IN1(n6254), .IN2(n5641), .IN3(n5646), .IN4(n2035), .Q(n2034)
         );
  OA22X1 U2303 ( .IN1(n5625), .IN2(n2036), .IN3(n6258), .IN4(n5633), .Q(n2035)
         );
  OA22X1 U2304 ( .IN1(n6100), .IN2(n5620), .IN3(n5623), .IN4(n2037), .Q(n2036)
         );
  OA22X1 U2305 ( .IN1(n5602), .IN2(n2038), .IN3(n6104), .IN4(n5611), .Q(n2037)
         );
  AOI22X1 U2306 ( .IN1(n5593), .IN2(\decodedPacket[1][80] ), .IN3(
        \decodedPacket[0][80] ), .IN4(n5589), .QN(n2038) );
  OAI22X1 U2307 ( .IN1(n5674), .IN2(n2039), .IN3(n6409), .IN4(n5680), .QN(
        N9749) );
  OA22X1 U2308 ( .IN1(n5656), .IN2(n2040), .IN3(n6411), .IN4(n5665), .Q(n2039)
         );
  OA22X1 U2309 ( .IN1(n6255), .IN2(n5641), .IN3(n5646), .IN4(n2041), .Q(n2040)
         );
  OA22X1 U2310 ( .IN1(n5625), .IN2(n2042), .IN3(n6257), .IN4(n5633), .Q(n2041)
         );
  OA22X1 U2311 ( .IN1(n6101), .IN2(n5620), .IN3(n5623), .IN4(n2043), .Q(n2042)
         );
  OA22X1 U2312 ( .IN1(n5602), .IN2(n2044), .IN3(n6103), .IN4(n5611), .Q(n2043)
         );
  AOI22X1 U2313 ( .IN1(n5593), .IN2(\decodedPacket[1][79] ), .IN3(
        \decodedPacket[0][79] ), .IN4(n5589), .QN(n2044) );
  OAI22X1 U2314 ( .IN1(n5674), .IN2(n2045), .IN3(n6401), .IN4(n5680), .QN(
        N9748) );
  OA22X1 U2315 ( .IN1(n5656), .IN2(n2046), .IN3(n6410), .IN4(n5665), .Q(n2045)
         );
  OA22X1 U2316 ( .IN1(n6247), .IN2(n5641), .IN3(n5646), .IN4(n2047), .Q(n2046)
         );
  OA22X1 U2317 ( .IN1(n5625), .IN2(n2048), .IN3(n6256), .IN4(n5633), .Q(n2047)
         );
  OA22X1 U2318 ( .IN1(n6093), .IN2(n5620), .IN3(n5623), .IN4(n2049), .Q(n2048)
         );
  OA22X1 U2319 ( .IN1(n5602), .IN2(n2050), .IN3(n6102), .IN4(n5611), .Q(n2049)
         );
  AOI22X1 U2320 ( .IN1(n5593), .IN2(\decodedPacket[1][78] ), .IN3(
        \decodedPacket[0][78] ), .IN4(n5589), .QN(n2050) );
  OAI22X1 U2321 ( .IN1(n5674), .IN2(n2051), .IN3(n6399), .IN4(n5678), .QN(
        N9747) );
  OA22X1 U2322 ( .IN1(n5656), .IN2(n2052), .IN3(n6352), .IN4(n5665), .Q(n2051)
         );
  OA22X1 U2323 ( .IN1(n6244), .IN2(n5641), .IN3(n5646), .IN4(n2053), .Q(n2052)
         );
  OA22X1 U2324 ( .IN1(n5625), .IN2(n2054), .IN3(n6198), .IN4(n5633), .Q(n2053)
         );
  OA22X1 U2325 ( .IN1(n6090), .IN2(n5620), .IN3(n5623), .IN4(n2055), .Q(n2054)
         );
  OA22X1 U2326 ( .IN1(n5603), .IN2(n2056), .IN3(n6044), .IN4(n5611), .Q(n2055)
         );
  AOI22X1 U2327 ( .IN1(n5593), .IN2(\decodedPacket[1][77] ), .IN3(
        \decodedPacket[0][77] ), .IN4(n5589), .QN(n2056) );
  OAI22X1 U2328 ( .IN1(n5674), .IN2(n2057), .IN3(n6398), .IN4(n5679), .QN(
        N9746) );
  OA22X1 U2329 ( .IN1(n5656), .IN2(n2058), .IN3(n6402), .IN4(n5665), .Q(n2057)
         );
  OA22X1 U2330 ( .IN1(n6243), .IN2(n5641), .IN3(n5646), .IN4(n2059), .Q(n2058)
         );
  OA22X1 U2331 ( .IN1(n5625), .IN2(n2060), .IN3(n6248), .IN4(n5633), .Q(n2059)
         );
  OA22X1 U2332 ( .IN1(n6089), .IN2(n5620), .IN3(n5623), .IN4(n2061), .Q(n2060)
         );
  OA22X1 U2333 ( .IN1(n5603), .IN2(n2062), .IN3(n6094), .IN4(n5611), .Q(n2061)
         );
  AOI22X1 U2334 ( .IN1(n5593), .IN2(\decodedPacket[1][76] ), .IN3(
        \decodedPacket[0][76] ), .IN4(n5589), .QN(n2062) );
  OAI22X1 U2335 ( .IN1(n5674), .IN2(n2063), .IN3(n6397), .IN4(n5677), .QN(
        N9745) );
  OA22X1 U2336 ( .IN1(n5656), .IN2(n2064), .IN3(n6403), .IN4(n5665), .Q(n2063)
         );
  OA22X1 U2337 ( .IN1(n6242), .IN2(n5641), .IN3(n5647), .IN4(n2065), .Q(n2064)
         );
  OA22X1 U2338 ( .IN1(n5625), .IN2(n2066), .IN3(n6249), .IN4(n5633), .Q(n2065)
         );
  OA22X1 U2339 ( .IN1(n6089), .IN2(n5620), .IN3(n5623), .IN4(n2067), .Q(n2066)
         );
  OA22X1 U2340 ( .IN1(n5603), .IN2(n2068), .IN3(n6095), .IN4(n5610), .Q(n2067)
         );
  AOI22X1 U2341 ( .IN1(n5594), .IN2(\decodedPacket[1][75] ), .IN3(
        \decodedPacket[0][75] ), .IN4(n5589), .QN(n2068) );
  OAI22X1 U2342 ( .IN1(n5674), .IN2(n2069), .IN3(n6396), .IN4(n5676), .QN(
        N9744) );
  OA22X1 U2343 ( .IN1(n5656), .IN2(n2070), .IN3(n6404), .IN4(n5666), .Q(n2069)
         );
  OA22X1 U2344 ( .IN1(n6241), .IN2(n5641), .IN3(n5647), .IN4(n2071), .Q(n2070)
         );
  OA22X1 U2345 ( .IN1(n5625), .IN2(n2072), .IN3(n6250), .IN4(n5633), .Q(n2071)
         );
  OA22X1 U2346 ( .IN1(n6088), .IN2(n5620), .IN3(n5623), .IN4(n2073), .Q(n2072)
         );
  OA22X1 U2347 ( .IN1(n5603), .IN2(n2074), .IN3(n6096), .IN4(n5610), .Q(n2073)
         );
  AOI22X1 U2348 ( .IN1(n5594), .IN2(\decodedPacket[1][74] ), .IN3(
        \decodedPacket[0][74] ), .IN4(n5589), .QN(n2074) );
  OAI22X1 U2349 ( .IN1(n5675), .IN2(n2075), .IN3(n6399), .IN4(n5681), .QN(
        N9743) );
  OA22X1 U2350 ( .IN1(n5657), .IN2(n2076), .IN3(n6405), .IN4(n5666), .Q(n2075)
         );
  OA22X1 U2351 ( .IN1(n6243), .IN2(n5641), .IN3(n5647), .IN4(n2077), .Q(n2076)
         );
  OA22X1 U2352 ( .IN1(n5625), .IN2(n2078), .IN3(n6251), .IN4(n5632), .Q(n2077)
         );
  OA22X1 U2353 ( .IN1(n6087), .IN2(n5620), .IN3(n5623), .IN4(n2079), .Q(n2078)
         );
  OA22X1 U2354 ( .IN1(n5603), .IN2(n2080), .IN3(n6097), .IN4(n5610), .Q(n2079)
         );
  AOI22X1 U2355 ( .IN1(n5594), .IN2(\decodedPacket[1][73] ), .IN3(
        \decodedPacket[0][73] ), .IN4(n5589), .QN(n2080) );
  OAI22X1 U2356 ( .IN1(n5675), .IN2(n2081), .IN3(n6394), .IN4(n5679), .QN(
        N9742) );
  OA22X1 U2357 ( .IN1(n5657), .IN2(n2082), .IN3(n6393), .IN4(n5666), .Q(n2081)
         );
  OA22X1 U2358 ( .IN1(n6240), .IN2(n5641), .IN3(n5647), .IN4(n2083), .Q(n2082)
         );
  OA22X1 U2359 ( .IN1(n5625), .IN2(n2084), .IN3(n6239), .IN4(n5632), .Q(n2083)
         );
  OA22X1 U2360 ( .IN1(n6086), .IN2(n5620), .IN3(n5623), .IN4(n2085), .Q(n2084)
         );
  OA22X1 U2361 ( .IN1(n5603), .IN2(n2086), .IN3(n6085), .IN4(n5610), .Q(n2085)
         );
  AOI22X1 U2362 ( .IN1(n5594), .IN2(\decodedPacket[1][72] ), .IN3(
        \decodedPacket[0][72] ), .IN4(n5589), .QN(n2086) );
  OAI22X1 U2363 ( .IN1(n5675), .IN2(n2087), .IN3(n6361), .IN4(n5679), .QN(
        N9741) );
  OA22X1 U2364 ( .IN1(n5657), .IN2(n2088), .IN3(n6360), .IN4(n5666), .Q(n2087)
         );
  OA22X1 U2365 ( .IN1(n6207), .IN2(n5641), .IN3(n5647), .IN4(n2089), .Q(n2088)
         );
  OA22X1 U2366 ( .IN1(n5625), .IN2(n2090), .IN3(n6206), .IN4(n5632), .Q(n2089)
         );
  OA22X1 U2367 ( .IN1(n6053), .IN2(n5620), .IN3(n5623), .IN4(n2091), .Q(n2090)
         );
  OA22X1 U2368 ( .IN1(n5603), .IN2(n2092), .IN3(n6052), .IN4(n5610), .Q(n2091)
         );
  AOI22X1 U2369 ( .IN1(n5594), .IN2(\decodedPacket[1][71] ), .IN3(
        \decodedPacket[0][71] ), .IN4(n5589), .QN(n2092) );
  OAI22X1 U2370 ( .IN1(n5675), .IN2(n2093), .IN3(n6350), .IN4(n5679), .QN(
        N9740) );
  OA22X1 U2371 ( .IN1(n5657), .IN2(n2094), .IN3(n6351), .IN4(n5666), .Q(n2093)
         );
  OA22X1 U2372 ( .IN1(n6196), .IN2(n5641), .IN3(n5644), .IN4(n2095), .Q(n2094)
         );
  OA22X1 U2373 ( .IN1(n5625), .IN2(n2096), .IN3(n6197), .IN4(n5632), .Q(n2095)
         );
  OA22X1 U2374 ( .IN1(n6042), .IN2(n5619), .IN3(n5623), .IN4(n2097), .Q(n2096)
         );
  OA22X1 U2375 ( .IN1(n5603), .IN2(n2098), .IN3(n6043), .IN4(n5609), .Q(n2097)
         );
  AOI22X1 U2376 ( .IN1(n5594), .IN2(\decodedPacket[1][70] ), .IN3(
        \decodedPacket[0][70] ), .IN4(n5590), .QN(n2098) );
  OAI22X1 U2377 ( .IN1(n5675), .IN2(n2099), .IN3(n6395), .IN4(n5679), .QN(
        N9739) );
  OA22X1 U2378 ( .IN1(n5657), .IN2(n2100), .IN3(n6392), .IN4(n5666), .Q(n2099)
         );
  OA22X1 U2379 ( .IN1(n6245), .IN2(n5640), .IN3(n5646), .IN4(n2101), .Q(n2100)
         );
  OA22X1 U2380 ( .IN1(n5625), .IN2(n2102), .IN3(n6238), .IN4(n5632), .Q(n2101)
         );
  OA22X1 U2381 ( .IN1(n6091), .IN2(n5619), .IN3(n5623), .IN4(n2103), .Q(n2102)
         );
  OA22X1 U2382 ( .IN1(n5603), .IN2(n2104), .IN3(n6084), .IN4(n5609), .Q(n2103)
         );
  AOI22X1 U2383 ( .IN1(n5594), .IN2(\decodedPacket[1][69] ), .IN3(
        \decodedPacket[0][69] ), .IN4(n5590), .QN(n2104) );
  OAI22X1 U2384 ( .IN1(n5675), .IN2(n2105), .IN3(n6423), .IN4(n5679), .QN(
        N9738) );
  OA22X1 U2385 ( .IN1(n5657), .IN2(n2106), .IN3(n6423), .IN4(n5666), .Q(n2105)
         );
  OA22X1 U2386 ( .IN1(n6269), .IN2(n5640), .IN3(n5649), .IN4(n2107), .Q(n2106)
         );
  OA22X1 U2387 ( .IN1(n5625), .IN2(n2108), .IN3(n6269), .IN4(n5632), .Q(n2107)
         );
  OA22X1 U2388 ( .IN1(n6115), .IN2(n5619), .IN3(n5622), .IN4(n2109), .Q(n2108)
         );
  OA22X1 U2389 ( .IN1(n5603), .IN2(n2110), .IN3(n6115), .IN4(n5609), .Q(n2109)
         );
  AOI22X1 U2390 ( .IN1(n5594), .IN2(\decodedPacket[1][68] ), .IN3(
        \decodedPacket[0][68] ), .IN4(n5590), .QN(n2110) );
  OAI22X1 U2391 ( .IN1(n5675), .IN2(n2111), .IN3(n6424), .IN4(n5679), .QN(
        N9737) );
  OA22X1 U2392 ( .IN1(n5657), .IN2(n2112), .IN3(n6424), .IN4(n5666), .Q(n2111)
         );
  OA22X1 U2393 ( .IN1(n6270), .IN2(n5640), .IN3(n5644), .IN4(n2113), .Q(n2112)
         );
  OA22X1 U2394 ( .IN1(n5625), .IN2(n2114), .IN3(n6270), .IN4(n5632), .Q(n2113)
         );
  OA22X1 U2395 ( .IN1(n6116), .IN2(n5619), .IN3(n5200), .IN4(n2115), .Q(n2114)
         );
  OA22X1 U2396 ( .IN1(n5603), .IN2(n2116), .IN3(n6116), .IN4(n5609), .Q(n2115)
         );
  AOI22X1 U2397 ( .IN1(n5594), .IN2(\decodedPacket[1][67] ), .IN3(
        \decodedPacket[0][67] ), .IN4(n5590), .QN(n2116) );
  OAI22X1 U2398 ( .IN1(n5675), .IN2(n2117), .IN3(n6425), .IN4(n5678), .QN(
        N9736) );
  OA22X1 U2399 ( .IN1(n5657), .IN2(n2118), .IN3(n6425), .IN4(n5666), .Q(n2117)
         );
  OA22X1 U2400 ( .IN1(n6271), .IN2(n5640), .IN3(n5645), .IN4(n2119), .Q(n2118)
         );
  OA22X1 U2401 ( .IN1(n5625), .IN2(n2120), .IN3(n6271), .IN4(n5632), .Q(n2119)
         );
  OA22X1 U2402 ( .IN1(n6117), .IN2(n5619), .IN3(n5200), .IN4(n2121), .Q(n2120)
         );
  OA22X1 U2403 ( .IN1(n5603), .IN2(n2122), .IN3(n6117), .IN4(n5609), .Q(n2121)
         );
  AOI22X1 U2404 ( .IN1(n5594), .IN2(\decodedPacket[1][66] ), .IN3(
        \decodedPacket[0][66] ), .IN4(n5590), .QN(n2122) );
  OAI22X1 U2405 ( .IN1(n5675), .IN2(n2123), .IN3(n6426), .IN4(n5678), .QN(
        N9735) );
  OA22X1 U2406 ( .IN1(n5657), .IN2(n2124), .IN3(n6426), .IN4(n5666), .Q(n2123)
         );
  OA22X1 U2407 ( .IN1(n6272), .IN2(n5640), .IN3(n5643), .IN4(n2125), .Q(n2124)
         );
  OA22X1 U2408 ( .IN1(n5625), .IN2(n2126), .IN3(n6272), .IN4(n5632), .Q(n2125)
         );
  OA22X1 U2409 ( .IN1(n6118), .IN2(n5619), .IN3(n5200), .IN4(n2127), .Q(n2126)
         );
  OA22X1 U2410 ( .IN1(n5603), .IN2(n2128), .IN3(n6118), .IN4(n5608), .Q(n2127)
         );
  AOI22X1 U2411 ( .IN1(n5594), .IN2(\decodedPacket[1][65] ), .IN3(
        \decodedPacket[0][65] ), .IN4(n5590), .QN(n2128) );
  OAI22X1 U2412 ( .IN1(n5675), .IN2(n2129), .IN3(n6427), .IN4(n5678), .QN(
        N9734) );
  OA22X1 U2413 ( .IN1(n5657), .IN2(n2130), .IN3(n6427), .IN4(n5666), .Q(n2129)
         );
  OA22X1 U2414 ( .IN1(n6273), .IN2(n5640), .IN3(n5648), .IN4(n2131), .Q(n2130)
         );
  OA22X1 U2415 ( .IN1(n5625), .IN2(n2132), .IN3(n6273), .IN4(n5632), .Q(n2131)
         );
  OA22X1 U2416 ( .IN1(n6119), .IN2(n5619), .IN3(n5200), .IN4(n2133), .Q(n2132)
         );
  OA22X1 U2417 ( .IN1(n5603), .IN2(n2134), .IN3(n6119), .IN4(n5608), .Q(n2133)
         );
  AOI22X1 U2418 ( .IN1(n5594), .IN2(\decodedPacket[1][64] ), .IN3(
        \decodedPacket[0][64] ), .IN4(n5590), .QN(n2134) );
  OAI22X1 U2419 ( .IN1(n5675), .IN2(n2135), .IN3(n6428), .IN4(n5678), .QN(
        N9733) );
  OA22X1 U2420 ( .IN1(n5657), .IN2(n2136), .IN3(n6428), .IN4(n5666), .Q(n2135)
         );
  OA22X1 U2421 ( .IN1(n6274), .IN2(n5640), .IN3(n5648), .IN4(n2137), .Q(n2136)
         );
  OA22X1 U2422 ( .IN1(n5625), .IN2(n2138), .IN3(n6274), .IN4(n5632), .Q(n2137)
         );
  OA22X1 U2423 ( .IN1(n6120), .IN2(n5619), .IN3(n5200), .IN4(n2139), .Q(n2138)
         );
  OA22X1 U2424 ( .IN1(n5603), .IN2(n2140), .IN3(n6120), .IN4(n5608), .Q(n2139)
         );
  AOI22X1 U2425 ( .IN1(n5594), .IN2(\decodedPacket[1][63] ), .IN3(
        \decodedPacket[0][63] ), .IN4(n5590), .QN(n2140) );
  OAI22X1 U2426 ( .IN1(n5675), .IN2(n2141), .IN3(n6429), .IN4(n5678), .QN(
        N9732) );
  OA22X1 U2427 ( .IN1(n5657), .IN2(n2142), .IN3(n6429), .IN4(n5666), .Q(n2141)
         );
  OA22X1 U2428 ( .IN1(n6275), .IN2(n5640), .IN3(n5643), .IN4(n2143), .Q(n2142)
         );
  OA22X1 U2429 ( .IN1(n5625), .IN2(n2144), .IN3(n6275), .IN4(n5632), .Q(n2143)
         );
  OA22X1 U2430 ( .IN1(n6121), .IN2(n5619), .IN3(n5200), .IN4(n2145), .Q(n2144)
         );
  OA22X1 U2431 ( .IN1(n5604), .IN2(n2146), .IN3(n6121), .IN4(n5608), .Q(n2145)
         );
  AOI22X1 U2432 ( .IN1(n5594), .IN2(\decodedPacket[1][62] ), .IN3(
        \decodedPacket[0][62] ), .IN4(n5590), .QN(n2146) );
  OAI22X1 U2433 ( .IN1(n5675), .IN2(n2147), .IN3(n6430), .IN4(n5678), .QN(
        N9731) );
  OA22X1 U2434 ( .IN1(n5658), .IN2(n2148), .IN3(n6430), .IN4(n5666), .Q(n2147)
         );
  OA22X1 U2435 ( .IN1(n6276), .IN2(n5640), .IN3(n5650), .IN4(n2149), .Q(n2148)
         );
  OA22X1 U2436 ( .IN1(n5625), .IN2(n2150), .IN3(n6276), .IN4(n5632), .Q(n2149)
         );
  OA22X1 U2437 ( .IN1(n6122), .IN2(n5619), .IN3(n5200), .IN4(n2151), .Q(n2150)
         );
  OA22X1 U2438 ( .IN1(n5604), .IN2(n2152), .IN3(n6122), .IN4(n5608), .Q(n2151)
         );
  AOI22X1 U2439 ( .IN1(n5594), .IN2(\decodedPacket[1][61] ), .IN3(
        \decodedPacket[0][61] ), .IN4(n5590), .QN(n2152) );
  OAI22X1 U2440 ( .IN1(n5675), .IN2(n2153), .IN3(n6431), .IN4(n5677), .QN(
        N9730) );
  OA22X1 U2441 ( .IN1(n5658), .IN2(n2154), .IN3(n6431), .IN4(n5667), .Q(n2153)
         );
  OA22X1 U2442 ( .IN1(n6277), .IN2(n5640), .IN3(n5648), .IN4(n2155), .Q(n2154)
         );
  OA22X1 U2443 ( .IN1(n5625), .IN2(n2156), .IN3(n6277), .IN4(n5631), .Q(n2155)
         );
  OA22X1 U2444 ( .IN1(n6123), .IN2(n5619), .IN3(n5200), .IN4(n2157), .Q(n2156)
         );
  OA22X1 U2445 ( .IN1(n5604), .IN2(n2158), .IN3(n6123), .IN4(n5597), .Q(n2157)
         );
  AOI22X1 U2446 ( .IN1(n5594), .IN2(\decodedPacket[1][60] ), .IN3(
        \decodedPacket[0][60] ), .IN4(n5590), .QN(n2158) );
  OAI22X1 U2447 ( .IN1(n5675), .IN2(n2159), .IN3(n6432), .IN4(n5677), .QN(
        N9729) );
  OA22X1 U2448 ( .IN1(n5658), .IN2(n2160), .IN3(n6432), .IN4(n5667), .Q(n2159)
         );
  OA22X1 U2449 ( .IN1(n6278), .IN2(n5640), .IN3(n5648), .IN4(n2161), .Q(n2160)
         );
  OA22X1 U2450 ( .IN1(n5625), .IN2(n2162), .IN3(n6278), .IN4(n5631), .Q(n2161)
         );
  OA22X1 U2451 ( .IN1(n6124), .IN2(n5619), .IN3(n5200), .IN4(n2163), .Q(n2162)
         );
  OA22X1 U2452 ( .IN1(n5604), .IN2(n2164), .IN3(n6124), .IN4(n5598), .Q(n2163)
         );
  AOI22X1 U2453 ( .IN1(n5594), .IN2(\decodedPacket[1][59] ), .IN3(
        \decodedPacket[0][59] ), .IN4(n5590), .QN(n2164) );
  OAI22X1 U2454 ( .IN1(n5675), .IN2(n2165), .IN3(n6433), .IN4(n5677), .QN(
        N9728) );
  OA22X1 U2455 ( .IN1(n5658), .IN2(n2166), .IN3(n6433), .IN4(n5667), .Q(n2165)
         );
  OA22X1 U2456 ( .IN1(n6279), .IN2(n5640), .IN3(n5648), .IN4(n2167), .Q(n2166)
         );
  OA22X1 U2457 ( .IN1(n5625), .IN2(n2168), .IN3(n6279), .IN4(n5631), .Q(n2167)
         );
  OA22X1 U2458 ( .IN1(n6125), .IN2(n5619), .IN3(n5622), .IN4(n2169), .Q(n2168)
         );
  OA22X1 U2459 ( .IN1(n5604), .IN2(n2170), .IN3(n6125), .IN4(n5599), .Q(n2169)
         );
  AOI22X1 U2460 ( .IN1(n5595), .IN2(\decodedPacket[1][58] ), .IN3(
        \decodedPacket[0][58] ), .IN4(n5590), .QN(n2170) );
  OAI22X1 U2461 ( .IN1(n5675), .IN2(n2171), .IN3(n6434), .IN4(n5677), .QN(
        N9727) );
  OA22X1 U2462 ( .IN1(n5658), .IN2(n2172), .IN3(n6434), .IN4(n5667), .Q(n2171)
         );
  OA22X1 U2463 ( .IN1(n6280), .IN2(n5640), .IN3(n5648), .IN4(n2173), .Q(n2172)
         );
  OA22X1 U2464 ( .IN1(n5625), .IN2(n2174), .IN3(n6280), .IN4(n5631), .Q(n2173)
         );
  OA22X1 U2465 ( .IN1(n6126), .IN2(n5619), .IN3(n5622), .IN4(n2175), .Q(n2174)
         );
  OA22X1 U2466 ( .IN1(n5604), .IN2(n2176), .IN3(n6126), .IN4(n5598), .Q(n2175)
         );
  AOI22X1 U2467 ( .IN1(n5595), .IN2(\decodedPacket[1][57] ), .IN3(
        \decodedPacket[0][57] ), .IN4(n5590), .QN(n2176) );
  OAI22X1 U2468 ( .IN1(n5675), .IN2(n2177), .IN3(n6435), .IN4(n5677), .QN(
        N9726) );
  OA22X1 U2469 ( .IN1(n5658), .IN2(n2178), .IN3(n6435), .IN4(n5667), .Q(n2177)
         );
  OA22X1 U2470 ( .IN1(n6281), .IN2(n5640), .IN3(n5648), .IN4(n2179), .Q(n2178)
         );
  OA22X1 U2471 ( .IN1(n5626), .IN2(n2180), .IN3(n6281), .IN4(n5631), .Q(n2179)
         );
  OA22X1 U2472 ( .IN1(n6127), .IN2(n5619), .IN3(n5622), .IN4(n2181), .Q(n2180)
         );
  OA22X1 U2473 ( .IN1(n5604), .IN2(n2182), .IN3(n6127), .IN4(n5610), .Q(n2181)
         );
  AOI22X1 U2474 ( .IN1(n5595), .IN2(\decodedPacket[1][56] ), .IN3(
        \decodedPacket[0][56] ), .IN4(n5590), .QN(n2182) );
  OAI22X1 U2475 ( .IN1(n5675), .IN2(n2183), .IN3(n6436), .IN4(n5677), .QN(
        N9725) );
  OA22X1 U2476 ( .IN1(n5658), .IN2(n2184), .IN3(n6436), .IN4(n5667), .Q(n2183)
         );
  OA22X1 U2477 ( .IN1(n6282), .IN2(n5640), .IN3(n5649), .IN4(n2185), .Q(n2184)
         );
  OA22X1 U2478 ( .IN1(n5626), .IN2(n2186), .IN3(n6282), .IN4(n5631), .Q(n2185)
         );
  OA22X1 U2479 ( .IN1(n6128), .IN2(n5619), .IN3(n5622), .IN4(n2187), .Q(n2186)
         );
  OA22X1 U2480 ( .IN1(n5604), .IN2(n2188), .IN3(n6128), .IN4(n5608), .Q(n2187)
         );
  AOI22X1 U2481 ( .IN1(n5595), .IN2(\decodedPacket[1][55] ), .IN3(
        \decodedPacket[0][55] ), .IN4(n5590), .QN(n2188) );
  OAI22X1 U2482 ( .IN1(n5675), .IN2(n2189), .IN3(n6437), .IN4(n5676), .QN(
        N9724) );
  OA22X1 U2483 ( .IN1(n5658), .IN2(n2190), .IN3(n6437), .IN4(n5667), .Q(n2189)
         );
  OA22X1 U2484 ( .IN1(n6283), .IN2(n5640), .IN3(n5649), .IN4(n2191), .Q(n2190)
         );
  OA22X1 U2485 ( .IN1(n5626), .IN2(n2192), .IN3(n6283), .IN4(n5631), .Q(n2191)
         );
  OA22X1 U2486 ( .IN1(n6129), .IN2(n5619), .IN3(n5622), .IN4(n2193), .Q(n2192)
         );
  OA22X1 U2487 ( .IN1(n5604), .IN2(n2194), .IN3(n6129), .IN4(n5609), .Q(n2193)
         );
  AOI22X1 U2488 ( .IN1(n5595), .IN2(\decodedPacket[1][54] ), .IN3(
        \decodedPacket[0][54] ), .IN4(n5590), .QN(n2194) );
  OAI22X1 U2489 ( .IN1(n5675), .IN2(n2195), .IN3(n6438), .IN4(n5676), .QN(
        N9723) );
  OA22X1 U2490 ( .IN1(n5658), .IN2(n2196), .IN3(n6438), .IN4(n5667), .Q(n2195)
         );
  OA22X1 U2491 ( .IN1(n6284), .IN2(n5640), .IN3(n5649), .IN4(n2197), .Q(n2196)
         );
  OA22X1 U2492 ( .IN1(n5626), .IN2(n2198), .IN3(n6284), .IN4(n5631), .Q(n2197)
         );
  OA22X1 U2493 ( .IN1(n6130), .IN2(n5619), .IN3(n5622), .IN4(n2199), .Q(n2198)
         );
  OA22X1 U2494 ( .IN1(n5604), .IN2(n2200), .IN3(n6130), .IN4(n5610), .Q(n2199)
         );
  AOI22X1 U2495 ( .IN1(n5595), .IN2(\decodedPacket[1][53] ), .IN3(
        \decodedPacket[0][53] ), .IN4(n5590), .QN(n2200) );
  OAI22X1 U2496 ( .IN1(n5675), .IN2(n2201), .IN3(n6439), .IN4(n5676), .QN(
        N9722) );
  OA22X1 U2497 ( .IN1(n5658), .IN2(n2202), .IN3(n6439), .IN4(n5667), .Q(n2201)
         );
  OA22X1 U2498 ( .IN1(n6285), .IN2(n5640), .IN3(n5649), .IN4(n2203), .Q(n2202)
         );
  OA22X1 U2499 ( .IN1(n5626), .IN2(n2204), .IN3(n6285), .IN4(n5631), .Q(n2203)
         );
  OA22X1 U2500 ( .IN1(n6131), .IN2(n5619), .IN3(n5622), .IN4(n2205), .Q(n2204)
         );
  OA22X1 U2501 ( .IN1(n5604), .IN2(n2206), .IN3(n6131), .IN4(n5611), .Q(n2205)
         );
  AOI22X1 U2502 ( .IN1(n5595), .IN2(\decodedPacket[1][52] ), .IN3(
        \decodedPacket[0][52] ), .IN4(n5590), .QN(n2206) );
  OAI22X1 U2503 ( .IN1(n5675), .IN2(n2207), .IN3(n6440), .IN4(n5676), .QN(
        N9721) );
  OA22X1 U2504 ( .IN1(n5658), .IN2(n2208), .IN3(n6440), .IN4(n5667), .Q(n2207)
         );
  OA22X1 U2505 ( .IN1(n6286), .IN2(n5640), .IN3(n5649), .IN4(n2209), .Q(n2208)
         );
  OA22X1 U2506 ( .IN1(n5626), .IN2(n2210), .IN3(n6286), .IN4(n5631), .Q(n2209)
         );
  OA22X1 U2507 ( .IN1(n6132), .IN2(n5619), .IN3(n5622), .IN4(n2211), .Q(n2210)
         );
  OA22X1 U2508 ( .IN1(n5604), .IN2(n2212), .IN3(n6132), .IN4(n5613), .Q(n2211)
         );
  AOI22X1 U2509 ( .IN1(n5595), .IN2(\decodedPacket[1][51] ), .IN3(
        \decodedPacket[0][51] ), .IN4(n5590), .QN(n2212) );
  OAI22X1 U2510 ( .IN1(n5675), .IN2(n2213), .IN3(n6441), .IN4(n5676), .QN(
        N9720) );
  OA22X1 U2511 ( .IN1(n5658), .IN2(n2214), .IN3(n6441), .IN4(n5667), .Q(n2213)
         );
  OA22X1 U2512 ( .IN1(n6287), .IN2(n5640), .IN3(n5650), .IN4(n2215), .Q(n2214)
         );
  OA22X1 U2513 ( .IN1(n5626), .IN2(n2216), .IN3(n6287), .IN4(n5631), .Q(n2215)
         );
  OA22X1 U2514 ( .IN1(n6133), .IN2(n5619), .IN3(n5622), .IN4(n2217), .Q(n2216)
         );
  OA22X1 U2515 ( .IN1(n5604), .IN2(n2218), .IN3(n6133), .IN4(n5611), .Q(n2217)
         );
  AOI22X1 U2516 ( .IN1(n5595), .IN2(\decodedPacket[1][50] ), .IN3(
        \decodedPacket[0][50] ), .IN4(n5590), .QN(n2218) );
  OAI22X1 U2517 ( .IN1(n5675), .IN2(n2219), .IN3(n6442), .IN4(n5676), .QN(
        N9719) );
  OA22X1 U2518 ( .IN1(n5659), .IN2(n2220), .IN3(n6442), .IN4(n5667), .Q(n2219)
         );
  OA22X1 U2519 ( .IN1(n6288), .IN2(n5640), .IN3(n5650), .IN4(n2221), .Q(n2220)
         );
  OA22X1 U2520 ( .IN1(n5626), .IN2(n2222), .IN3(n6288), .IN4(n5631), .Q(n2221)
         );
  OA22X1 U2521 ( .IN1(n6134), .IN2(n5619), .IN3(n5622), .IN4(n2223), .Q(n2222)
         );
  OA22X1 U2522 ( .IN1(n5604), .IN2(n2224), .IN3(n6134), .IN4(n5613), .Q(n2223)
         );
  AOI22X1 U2523 ( .IN1(n5595), .IN2(\decodedPacket[1][49] ), .IN3(
        \decodedPacket[0][49] ), .IN4(n5590), .QN(n2224) );
  OAI22X1 U2524 ( .IN1(n5675), .IN2(n2225), .IN3(n6443), .IN4(n5682), .QN(
        N9718) );
  OA22X1 U2525 ( .IN1(n5659), .IN2(n2226), .IN3(n6443), .IN4(n5667), .Q(n2225)
         );
  OA22X1 U2526 ( .IN1(n6289), .IN2(n5640), .IN3(n5650), .IN4(n2227), .Q(n2226)
         );
  OA22X1 U2527 ( .IN1(n5626), .IN2(n2228), .IN3(n6289), .IN4(n5631), .Q(n2227)
         );
  OA22X1 U2528 ( .IN1(n6135), .IN2(n5619), .IN3(n5622), .IN4(n2229), .Q(n2228)
         );
  OA22X1 U2529 ( .IN1(n5604), .IN2(n2230), .IN3(n6135), .IN4(n5611), .Q(n2229)
         );
  AOI22X1 U2530 ( .IN1(n5595), .IN2(\decodedPacket[1][48] ), .IN3(
        \decodedPacket[0][48] ), .IN4(n5590), .QN(n2230) );
  OAI22X1 U2531 ( .IN1(n5675), .IN2(n2231), .IN3(n6444), .IN4(n5680), .QN(
        N9716) );
  OA22X1 U2532 ( .IN1(n5659), .IN2(n2232), .IN3(n6444), .IN4(n5667), .Q(n2231)
         );
  OA22X1 U2533 ( .IN1(n6290), .IN2(n5640), .IN3(n5650), .IN4(n2233), .Q(n2232)
         );
  OA22X1 U2534 ( .IN1(n5626), .IN2(n2234), .IN3(n6290), .IN4(n5630), .Q(n2233)
         );
  OA22X1 U2535 ( .IN1(n6136), .IN2(n5619), .IN3(n5622), .IN4(n2235), .Q(n2234)
         );
  OA22X1 U2536 ( .IN1(n5605), .IN2(n2236), .IN3(n6136), .IN4(n5597), .Q(n2235)
         );
  AOI22X1 U2537 ( .IN1(n5595), .IN2(\decodedPacket[1][47] ), .IN3(
        \decodedPacket[0][47] ), .IN4(n5590), .QN(n2236) );
  OAI22X1 U2538 ( .IN1(n5675), .IN2(n2237), .IN3(n6445), .IN4(n5678), .QN(
        N9715) );
  OA22X1 U2539 ( .IN1(n5659), .IN2(n2238), .IN3(n6445), .IN4(n5667), .Q(n2237)
         );
  OA22X1 U2540 ( .IN1(n6291), .IN2(n5640), .IN3(n5650), .IN4(n2239), .Q(n2238)
         );
  OA22X1 U2541 ( .IN1(n5626), .IN2(n2240), .IN3(n6291), .IN4(n5630), .Q(n2239)
         );
  OA22X1 U2542 ( .IN1(n6137), .IN2(n5619), .IN3(n5622), .IN4(n2241), .Q(n2240)
         );
  OA22X1 U2543 ( .IN1(n5605), .IN2(n2242), .IN3(n6137), .IN4(n5598), .Q(n2241)
         );
  AOI22X1 U2544 ( .IN1(n5595), .IN2(\decodedPacket[1][46] ), .IN3(
        \decodedPacket[0][46] ), .IN4(n5590), .QN(n2242) );
  OAI22X1 U2545 ( .IN1(n5675), .IN2(n2243), .IN3(n6446), .IN4(n5677), .QN(
        N9714) );
  OA22X1 U2546 ( .IN1(n5659), .IN2(n2244), .IN3(n6446), .IN4(n5668), .Q(n2243)
         );
  OA22X1 U2547 ( .IN1(n6292), .IN2(n5640), .IN3(n5646), .IN4(n2245), .Q(n2244)
         );
  OA22X1 U2548 ( .IN1(n5626), .IN2(n2246), .IN3(n6292), .IN4(n5630), .Q(n2245)
         );
  OA22X1 U2549 ( .IN1(n6138), .IN2(n5619), .IN3(n5622), .IN4(n2247), .Q(n2246)
         );
  OA22X1 U2550 ( .IN1(n5605), .IN2(n2248), .IN3(n6138), .IN4(n5615), .Q(n2247)
         );
  AOI22X1 U2551 ( .IN1(n5595), .IN2(\decodedPacket[1][45] ), .IN3(
        \decodedPacket[0][45] ), .IN4(n5590), .QN(n2248) );
  OAI22X1 U2552 ( .IN1(n5675), .IN2(n2249), .IN3(n6447), .IN4(n5676), .QN(
        N9713) );
  OA22X1 U2553 ( .IN1(n5659), .IN2(n2250), .IN3(n6447), .IN4(n5668), .Q(n2249)
         );
  OA22X1 U2554 ( .IN1(n6293), .IN2(n5640), .IN3(n5650), .IN4(n2251), .Q(n2250)
         );
  OA22X1 U2555 ( .IN1(n5626), .IN2(n2252), .IN3(n6293), .IN4(n5630), .Q(n2251)
         );
  OA22X1 U2556 ( .IN1(n6139), .IN2(n5619), .IN3(n5622), .IN4(n2253), .Q(n2252)
         );
  OA22X1 U2557 ( .IN1(n5605), .IN2(n2254), .IN3(n6139), .IN4(n5608), .Q(n2253)
         );
  AOI22X1 U2558 ( .IN1(n5595), .IN2(\decodedPacket[1][44] ), .IN3(
        \decodedPacket[0][44] ), .IN4(n5590), .QN(n2254) );
  OAI22X1 U2559 ( .IN1(n5675), .IN2(n2255), .IN3(n6448), .IN4(n5681), .QN(
        N9712) );
  OA22X1 U2560 ( .IN1(n5659), .IN2(n2256), .IN3(n6448), .IN4(n5668), .Q(n2255)
         );
  OA22X1 U2561 ( .IN1(n6294), .IN2(n5640), .IN3(n5647), .IN4(n2257), .Q(n2256)
         );
  OA22X1 U2562 ( .IN1(n5626), .IN2(n2258), .IN3(n6294), .IN4(n5630), .Q(n2257)
         );
  OA22X1 U2563 ( .IN1(n6140), .IN2(n5619), .IN3(n5622), .IN4(n2259), .Q(n2258)
         );
  OA22X1 U2564 ( .IN1(n5605), .IN2(n2260), .IN3(n6140), .IN4(n5614), .Q(n2259)
         );
  AOI22X1 U2565 ( .IN1(n5595), .IN2(\decodedPacket[1][43] ), .IN3(
        \decodedPacket[0][43] ), .IN4(n5590), .QN(n2260) );
  OAI22X1 U2566 ( .IN1(n5675), .IN2(n2261), .IN3(n6449), .IN4(n5677), .QN(
        N9711) );
  OA22X1 U2567 ( .IN1(n5659), .IN2(n2262), .IN3(n6449), .IN4(n5668), .Q(n2261)
         );
  OA22X1 U2568 ( .IN1(n6295), .IN2(n5640), .IN3(n5648), .IN4(n2263), .Q(n2262)
         );
  OA22X1 U2569 ( .IN1(n5626), .IN2(n2264), .IN3(n6295), .IN4(n5630), .Q(n2263)
         );
  OA22X1 U2570 ( .IN1(n6141), .IN2(n5619), .IN3(n5622), .IN4(n2265), .Q(n2264)
         );
  OA22X1 U2571 ( .IN1(n5605), .IN2(n2266), .IN3(n6141), .IN4(n5608), .Q(n2265)
         );
  AOI22X1 U2572 ( .IN1(n5595), .IN2(\decodedPacket[1][42] ), .IN3(
        \decodedPacket[0][42] ), .IN4(n5590), .QN(n2266) );
  OAI22X1 U2573 ( .IN1(n5675), .IN2(n2267), .IN3(n6450), .IN4(n5676), .QN(
        N9710) );
  OA22X1 U2574 ( .IN1(n5659), .IN2(n2268), .IN3(n6450), .IN4(n5668), .Q(n2267)
         );
  OA22X1 U2575 ( .IN1(n6296), .IN2(n5640), .IN3(n5643), .IN4(n2269), .Q(n2268)
         );
  OA22X1 U2576 ( .IN1(n5626), .IN2(n2270), .IN3(n6296), .IN4(n5630), .Q(n2269)
         );
  OA22X1 U2577 ( .IN1(n6142), .IN2(n5619), .IN3(n5622), .IN4(n2271), .Q(n2270)
         );
  OA22X1 U2578 ( .IN1(n5605), .IN2(n2272), .IN3(n6142), .IN4(n5609), .Q(n2271)
         );
  AOI22X1 U2579 ( .IN1(n5596), .IN2(\decodedPacket[1][41] ), .IN3(
        \decodedPacket[0][41] ), .IN4(n5590), .QN(n2272) );
  OAI22X1 U2580 ( .IN1(n5675), .IN2(n2273), .IN3(n6451), .IN4(n5677), .QN(
        N9709) );
  OA22X1 U2581 ( .IN1(n5659), .IN2(n2274), .IN3(n6451), .IN4(n5668), .Q(n2273)
         );
  OA22X1 U2582 ( .IN1(n6297), .IN2(n5640), .IN3(n5645), .IN4(n2275), .Q(n2274)
         );
  OA22X1 U2583 ( .IN1(n5626), .IN2(n2276), .IN3(n6297), .IN4(n5630), .Q(n2275)
         );
  OA22X1 U2584 ( .IN1(n6143), .IN2(n5619), .IN3(n5622), .IN4(n2277), .Q(n2276)
         );
  OA22X1 U2585 ( .IN1(n5605), .IN2(n2278), .IN3(n6143), .IN4(n5613), .Q(n2277)
         );
  AOI22X1 U2586 ( .IN1(n5596), .IN2(\decodedPacket[1][40] ), .IN3(
        \decodedPacket[0][40] ), .IN4(n5590), .QN(n2278) );
  OAI22X1 U2587 ( .IN1(n5675), .IN2(n2279), .IN3(n6452), .IN4(n5682), .QN(
        N9708) );
  OA22X1 U2588 ( .IN1(n5659), .IN2(n2280), .IN3(n6452), .IN4(n5668), .Q(n2279)
         );
  OA22X1 U2589 ( .IN1(n6298), .IN2(n5640), .IN3(n5649), .IN4(n2281), .Q(n2280)
         );
  OA22X1 U2590 ( .IN1(n5626), .IN2(n2282), .IN3(n6298), .IN4(n5630), .Q(n2281)
         );
  OA22X1 U2591 ( .IN1(n6144), .IN2(n5619), .IN3(n5622), .IN4(n2283), .Q(n2282)
         );
  OA22X1 U2592 ( .IN1(n5605), .IN2(n2284), .IN3(n6144), .IN4(n5612), .Q(n2283)
         );
  AOI22X1 U2593 ( .IN1(n5596), .IN2(\decodedPacket[1][39] ), .IN3(
        \decodedPacket[0][39] ), .IN4(n5590), .QN(n2284) );
  OAI22X1 U2594 ( .IN1(n5675), .IN2(n2285), .IN3(n6453), .IN4(n5680), .QN(
        N9707) );
  OA22X1 U2595 ( .IN1(n5659), .IN2(n2286), .IN3(n6453), .IN4(n5668), .Q(n2285)
         );
  OA22X1 U2596 ( .IN1(n6299), .IN2(n5640), .IN3(n5646), .IN4(n2287), .Q(n2286)
         );
  OA22X1 U2597 ( .IN1(n5626), .IN2(n2288), .IN3(n6299), .IN4(n5630), .Q(n2287)
         );
  OA22X1 U2598 ( .IN1(n6145), .IN2(n5619), .IN3(n5622), .IN4(n2289), .Q(n2288)
         );
  OA22X1 U2599 ( .IN1(n5605), .IN2(n2290), .IN3(n6145), .IN4(n5608), .Q(n2289)
         );
  AOI22X1 U2600 ( .IN1(n5596), .IN2(\decodedPacket[1][38] ), .IN3(
        \decodedPacket[0][38] ), .IN4(n5590), .QN(n2290) );
  OAI22X1 U2601 ( .IN1(n5675), .IN2(n2291), .IN3(n6454), .IN4(n5678), .QN(
        N9706) );
  OA22X1 U2602 ( .IN1(n5660), .IN2(n2292), .IN3(n6454), .IN4(n5668), .Q(n2291)
         );
  OA22X1 U2603 ( .IN1(n6300), .IN2(n5640), .IN3(n5650), .IN4(n2293), .Q(n2292)
         );
  OA22X1 U2604 ( .IN1(n5626), .IN2(n2294), .IN3(n6300), .IN4(n5630), .Q(n2293)
         );
  OA22X1 U2605 ( .IN1(n6146), .IN2(n5618), .IN3(n5622), .IN4(n2295), .Q(n2294)
         );
  OA22X1 U2606 ( .IN1(n5605), .IN2(n2296), .IN3(n6146), .IN4(n5598), .Q(n2295)
         );
  AOI22X1 U2607 ( .IN1(n5596), .IN2(\decodedPacket[1][37] ), .IN3(
        \decodedPacket[0][37] ), .IN4(n5590), .QN(n2296) );
  OA22X1 U2609 ( .IN1(n5660), .IN2(n2298), .IN3(n6320), .IN4(n5668), .Q(n2297)
         );
  OA22X1 U2616 ( .IN1(n5660), .IN2(n2304), .IN3(n6321), .IN4(n5668), .Q(n2303)
         );
  OA22X1 U2623 ( .IN1(n5660), .IN2(n2310), .IN3(n6322), .IN4(n5668), .Q(n2309)
         );
  OA22X1 U2630 ( .IN1(n5660), .IN2(n2316), .IN3(n6323), .IN4(n5668), .Q(n2315)
         );
  OA22X1 U2637 ( .IN1(n5660), .IN2(n2322), .IN3(n6324), .IN4(n5668), .Q(n2321)
         );
  OA22X1 U2644 ( .IN1(n5660), .IN2(n2328), .IN3(n6325), .IN4(n5668), .Q(n2327)
         );
  OA22X1 U2651 ( .IN1(n5660), .IN2(n2334), .IN3(n6326), .IN4(n5669), .Q(n2333)
         );
  OA22X1 U2658 ( .IN1(n5660), .IN2(n2340), .IN3(n6327), .IN4(n5669), .Q(n2339)
         );
  OA22X1 U2665 ( .IN1(n5660), .IN2(n2346), .IN3(n6328), .IN4(n5669), .Q(n2345)
         );
  OA22X1 U2672 ( .IN1(n5660), .IN2(n2352), .IN3(n6329), .IN4(n5669), .Q(n2351)
         );
  OA22X1 U2679 ( .IN1(n5660), .IN2(n2358), .IN3(n6330), .IN4(n5669), .Q(n2357)
         );
  OA22X1 U2686 ( .IN1(n5661), .IN2(n2364), .IN3(n6331), .IN4(n5669), .Q(n2363)
         );
  OA22X1 U2693 ( .IN1(n5661), .IN2(n2370), .IN3(n6332), .IN4(n5669), .Q(n2369)
         );
  OA22X1 U2700 ( .IN1(n5661), .IN2(n2376), .IN3(n6333), .IN4(n5669), .Q(n2375)
         );
  OA22X1 U2707 ( .IN1(n5661), .IN2(n2382), .IN3(n6334), .IN4(n5669), .Q(n2381)
         );
  OA22X1 U2714 ( .IN1(n5661), .IN2(n2388), .IN3(n6335), .IN4(n5669), .Q(n2387)
         );
  OA22X1 U2721 ( .IN1(n5661), .IN2(n2394), .IN3(n6336), .IN4(n5669), .Q(n2393)
         );
  OA22X1 U2728 ( .IN1(n5661), .IN2(n2400), .IN3(n6337), .IN4(n5669), .Q(n2399)
         );
  OA22X1 U2735 ( .IN1(n5661), .IN2(n2406), .IN3(n6338), .IN4(n5669), .Q(n2405)
         );
  OA22X1 U2742 ( .IN1(n5661), .IN2(n2412), .IN3(n6339), .IN4(n5669), .Q(n2411)
         );
  OA22X1 U2749 ( .IN1(n5661), .IN2(n2418), .IN3(n6340), .IN4(n5669), .Q(n2417)
         );
  OA22X1 U2756 ( .IN1(n5661), .IN2(n2424), .IN3(n6341), .IN4(n5670), .Q(n2423)
         );
  OA22X1 U2763 ( .IN1(n5661), .IN2(n2430), .IN3(n6342), .IN4(n5670), .Q(n2429)
         );
  OA22X1 U2770 ( .IN1(n5662), .IN2(n2436), .IN3(n6343), .IN4(n5670), .Q(n2435)
         );
  OA22X1 U2777 ( .IN1(n5662), .IN2(n2442), .IN3(n6344), .IN4(n5670), .Q(n2441)
         );
  OA22X1 U2784 ( .IN1(n5662), .IN2(n2448), .IN3(n6345), .IN4(n5670), .Q(n2447)
         );
  OA22X1 U2791 ( .IN1(n5662), .IN2(n2454), .IN3(n6346), .IN4(n5670), .Q(n2453)
         );
  OA22X1 U2798 ( .IN1(n5662), .IN2(n2460), .IN3(n6315), .IN4(n5670), .Q(n2459)
         );
  OA22X1 U2805 ( .IN1(n5662), .IN2(n2466), .IN3(n6316), .IN4(n5670), .Q(n2465)
         );
  OA22X1 U2812 ( .IN1(n5662), .IN2(n2472), .IN3(n6317), .IN4(n5670), .Q(n2471)
         );
  OA22X1 U2819 ( .IN1(n5662), .IN2(n2478), .IN3(n6318), .IN4(n5670), .Q(n2477)
         );
  OA22X1 U2826 ( .IN1(n5662), .IN2(n2484), .IN3(n6319), .IN4(n5670), .Q(n2483)
         );
  OAI22X1 U2832 ( .IN1(n5675), .IN2(n2489), .IN3(n6455), .IN4(n5676), .QN(
        N9673) );
  OA22X1 U2833 ( .IN1(n5662), .IN2(n2490), .IN3(n6455), .IN4(n5670), .Q(n2489)
         );
  OA22X1 U2834 ( .IN1(n6301), .IN2(n5639), .IN3(n5647), .IN4(n2491), .Q(n2490)
         );
  OA22X1 U2835 ( .IN1(n5627), .IN2(n2492), .IN3(n6301), .IN4(n5636), .Q(n2491)
         );
  OA22X1 U2836 ( .IN1(n6147), .IN2(n5618), .IN3(n5622), .IN4(n2493), .Q(n2492)
         );
  OA22X1 U2837 ( .IN1(n5607), .IN2(n2494), .IN3(n6147), .IN4(n5611), .Q(n2493)
         );
  AOI22X1 U2838 ( .IN1(n5596), .IN2(\decodedPacket[1][4] ), .IN3(
        \decodedPacket[0][4] ), .IN4(n5590), .QN(n2494) );
  OAI22X1 U2839 ( .IN1(n5675), .IN2(n2495), .IN3(n6456), .IN4(n5677), .QN(
        N9672) );
  OA22X1 U2840 ( .IN1(n5662), .IN2(n2496), .IN3(n6456), .IN4(n5670), .Q(n2495)
         );
  OA22X1 U2841 ( .IN1(n6302), .IN2(n5639), .IN3(n5650), .IN4(n2497), .Q(n2496)
         );
  OA22X1 U2842 ( .IN1(n5627), .IN2(n2498), .IN3(n6302), .IN4(n5629), .Q(n2497)
         );
  OA22X1 U2843 ( .IN1(n6148), .IN2(n5618), .IN3(n5622), .IN4(n2499), .Q(n2498)
         );
  OA22X1 U2844 ( .IN1(n5607), .IN2(n2500), .IN3(n6148), .IN4(n5598), .Q(n2499)
         );
  AOI22X1 U2845 ( .IN1(n5596), .IN2(\decodedPacket[1][3] ), .IN3(
        \decodedPacket[0][3] ), .IN4(n5590), .QN(n2500) );
  OAI22X1 U2846 ( .IN1(n5675), .IN2(n2501), .IN3(n6457), .IN4(n5682), .QN(
        N9671) );
  OA22X1 U2847 ( .IN1(n5662), .IN2(n2502), .IN3(n6457), .IN4(n5670), .Q(n2501)
         );
  OA22X1 U2848 ( .IN1(n6303), .IN2(n5639), .IN3(n5647), .IN4(n2503), .Q(n2502)
         );
  OA22X1 U2849 ( .IN1(n5627), .IN2(n2504), .IN3(n6303), .IN4(n5628), .Q(n2503)
         );
  OA22X1 U2850 ( .IN1(n6149), .IN2(n5618), .IN3(n5622), .IN4(n2505), .Q(n2504)
         );
  OA22X1 U2851 ( .IN1(n5606), .IN2(n2506), .IN3(n6149), .IN4(n5612), .Q(n2505)
         );
  AOI22X1 U2852 ( .IN1(n5596), .IN2(\decodedPacket[1][2] ), .IN3(
        \decodedPacket[0][2] ), .IN4(n5590), .QN(n2506) );
  OAI22X1 U2853 ( .IN1(n5672), .IN2(n2507), .IN3(n6458), .IN4(n5680), .QN(
        N9670) );
  OA22X1 U2854 ( .IN1(n5654), .IN2(n2508), .IN3(n6458), .IN4(n5670), .Q(n2507)
         );
  OA22X1 U2855 ( .IN1(n6304), .IN2(n5639), .IN3(n5645), .IN4(n2509), .Q(n2508)
         );
  OA22X1 U2856 ( .IN1(n5627), .IN2(n2510), .IN3(n6304), .IN4(n5630), .Q(n2509)
         );
  OA22X1 U2857 ( .IN1(n6150), .IN2(n5618), .IN3(n5622), .IN4(n2511), .Q(n2510)
         );
  OA22X1 U2858 ( .IN1(n5607), .IN2(n2512), .IN3(n6150), .IN4(n5599), .Q(n2511)
         );
  AOI22X1 U2859 ( .IN1(n5596), .IN2(\decodedPacket[1][1] ), .IN3(
        \decodedPacket[0][1] ), .IN4(n5590), .QN(n2512) );
  OAI22X1 U2860 ( .IN1(n5671), .IN2(n2513), .IN3(n6459), .IN4(n5678), .QN(
        N9669) );
  OA22X1 U2861 ( .IN1(n5653), .IN2(n2514), .IN3(n6459), .IN4(n5663), .Q(n2513)
         );
  OA22X1 U2862 ( .IN1(n6305), .IN2(n5639), .IN3(n5649), .IN4(n2515), .Q(n2514)
         );
  OA22X1 U2863 ( .IN1(n5627), .IN2(n2516), .IN3(n6305), .IN4(n5636), .Q(n2515)
         );
  OA22X1 U2864 ( .IN1(n6151), .IN2(n5618), .IN3(n5623), .IN4(n2517), .Q(n2516)
         );
  OA22X1 U2865 ( .IN1(n5606), .IN2(n2518), .IN3(n6151), .IN4(n5613), .Q(n2517)
         );
  AOI22X1 U2866 ( .IN1(n5596), .IN2(\decodedPacket[1][0] ), .IN3(
        \decodedPacket[0][0] ), .IN4(n5590), .QN(n2518) );
  NAND4X0 U2867 ( .IN1(n5663), .IN2(n5639), .IN3(n2519), .IN4(n2520), .QN(
        decodedVector_o[0]) );
  NAND4X0 U2869 ( .IN1(n1752), .IN2(decodedPacketValid[7]), .IN3(n5992), .IN4(
        n5987), .QN(n1757) );
  NAND4X0 U2870 ( .IN1(n1754), .IN2(decodedPacketValid[4]), .IN3(n5995), .IN4(
        n5990), .QN(n1763) );
  NAND4X0 U2873 ( .IN1(n1753), .IN2(decodedPacketValid[6]), .IN3(n5993), .IN4(
        n5988), .QN(n1759) );
  OA21X1 U2875 ( .IN1(n5997), .IN2(decodedPacketValid[1]), .IN3(n5590), .Q(
        n2521) );
  OA22X1 U2893 ( .IN1(n5856), .IN2(n5561), .IN3(n5565), .IN4(n2540), .Q(n2539)
         );
  OAI22X1 U2896 ( .IN1(n6384), .IN2(n5585), .IN3(n5578), .IN4(n2542), .QN(
        N10701) );
  OA22X1 U2897 ( .IN1(n6349), .IN2(n5561), .IN3(n5571), .IN4(n2543), .Q(n2542)
         );
  OA22X1 U2898 ( .IN1(n5552), .IN2(n2544), .IN3(n6230), .IN4(n5544), .Q(n2543)
         );
  OA22X1 U2899 ( .IN1(n6195), .IN2(n5532), .IN3(n5275), .IN4(n6076), .Q(n2544)
         );
  OAI22X1 U2900 ( .IN1(n6376), .IN2(n5585), .IN3(n5578), .IN4(n2545), .QN(
        N10700) );
  OA22X1 U2901 ( .IN1(n6348), .IN2(n5561), .IN3(n5565), .IN4(n2546), .Q(n2545)
         );
  OA22X1 U2902 ( .IN1(n5552), .IN2(n2547), .IN3(n6222), .IN4(n5544), .Q(n2546)
         );
  OA22X1 U2903 ( .IN1(n6194), .IN2(n5532), .IN3(n5531), .IN4(n6068), .Q(n2547)
         );
  OAI22X1 U2904 ( .IN1(n6373), .IN2(n5585), .IN3(n5578), .IN4(n2548), .QN(
        N10699) );
  OA22X1 U2905 ( .IN1(n6374), .IN2(n5561), .IN3(n5562), .IN4(n2549), .Q(n2548)
         );
  OA22X1 U2906 ( .IN1(n5552), .IN2(n2550), .IN3(n6218), .IN4(n5544), .Q(n2549)
         );
  OA22X1 U2907 ( .IN1(n6220), .IN2(n5532), .IN3(n5531), .IN4(n6064), .Q(n2550)
         );
  OA22X1 U2909 ( .IN1(n6371), .IN2(n5561), .IN3(n5569), .IN4(n2552), .Q(n2551)
         );
  OAI22X1 U2912 ( .IN1(n6373), .IN2(n5585), .IN3(n5578), .IN4(n2554), .QN(
        N10697) );
  OA22X1 U2913 ( .IN1(n6370), .IN2(n5561), .IN3(n5568), .IN4(n2555), .Q(n2554)
         );
  OA22X1 U2914 ( .IN1(n5552), .IN2(n2556), .IN3(n6219), .IN4(n5544), .Q(n2555)
         );
  OA22X1 U2915 ( .IN1(n6216), .IN2(n5532), .IN3(n5531), .IN4(n6065), .Q(n2556)
         );
  OAI22X1 U2916 ( .IN1(n6397), .IN2(n5585), .IN3(n5579), .IN4(n2557), .QN(
        N10696) );
  OA22X1 U2917 ( .IN1(n6347), .IN2(n5561), .IN3(n5567), .IN4(n2558), .Q(n2557)
         );
  OA22X1 U2918 ( .IN1(n5551), .IN2(n2559), .IN3(n6245), .IN4(n5544), .Q(n2558)
         );
  OA22X1 U2919 ( .IN1(n6193), .IN2(n5532), .IN3(n5531), .IN4(n6091), .Q(n2559)
         );
  OAI22X1 U2920 ( .IN1(n5967), .IN2(n5585), .IN3(n5579), .IN4(n2560), .QN(
        N10695) );
  OA22X1 U2921 ( .IN1(n6369), .IN2(n5561), .IN3(n5562), .IN4(n2561), .Q(n2560)
         );
  OA22X1 U2922 ( .IN1(n5551), .IN2(n2562), .IN3(n5952), .IN4(n5544), .Q(n2561)
         );
  OA22X1 U2923 ( .IN1(n6215), .IN2(n5533), .IN3(n5531), .IN4(n5937), .Q(n2562)
         );
  OAI22X1 U2924 ( .IN1(n5968), .IN2(n5584), .IN3(n5579), .IN4(n2563), .QN(
        N10694) );
  OA22X1 U2925 ( .IN1(n6368), .IN2(n5561), .IN3(n5563), .IN4(n2564), .Q(n2563)
         );
  OA22X1 U2926 ( .IN1(n5551), .IN2(n2565), .IN3(n5953), .IN4(n5544), .Q(n2564)
         );
  OA22X1 U2927 ( .IN1(n6214), .IN2(n5533), .IN3(n5531), .IN4(n5938), .Q(n2565)
         );
  OAI22X1 U2928 ( .IN1(n5969), .IN2(n5584), .IN3(n5579), .IN4(n2566), .QN(
        N10693) );
  OA22X1 U2929 ( .IN1(n6367), .IN2(n5561), .IN3(n5564), .IN4(n2567), .Q(n2566)
         );
  OA22X1 U2930 ( .IN1(n5551), .IN2(n2568), .IN3(n5954), .IN4(n5544), .Q(n2567)
         );
  OA22X1 U2931 ( .IN1(n6213), .IN2(n5533), .IN3(n5531), .IN4(n5939), .Q(n2568)
         );
  OAI22X1 U2932 ( .IN1(n5970), .IN2(n5584), .IN3(n5579), .IN4(n2569), .QN(
        N10692) );
  OA22X1 U2933 ( .IN1(n6366), .IN2(n5561), .IN3(n5572), .IN4(n2570), .Q(n2569)
         );
  OA22X1 U2934 ( .IN1(n5551), .IN2(n2571), .IN3(n5955), .IN4(n5544), .Q(n2570)
         );
  OA22X1 U2935 ( .IN1(n6212), .IN2(n5533), .IN3(n5531), .IN4(n5940), .Q(n2571)
         );
  OAI22X1 U2936 ( .IN1(n5971), .IN2(n5584), .IN3(n5579), .IN4(n2572), .QN(
        N10691) );
  OA22X1 U2937 ( .IN1(n6365), .IN2(n5560), .IN3(n5566), .IN4(n2573), .Q(n2572)
         );
  OA22X1 U2938 ( .IN1(n5551), .IN2(n2574), .IN3(n5956), .IN4(n5544), .Q(n2573)
         );
  OA22X1 U2939 ( .IN1(n6211), .IN2(n5533), .IN3(n5531), .IN4(n5941), .Q(n2574)
         );
  OAI22X1 U2940 ( .IN1(n5972), .IN2(n5584), .IN3(n5579), .IN4(n2575), .QN(
        N10690) );
  OA22X1 U2941 ( .IN1(n6364), .IN2(n5560), .IN3(n5569), .IN4(n2576), .Q(n2575)
         );
  OA22X1 U2942 ( .IN1(n5551), .IN2(n2577), .IN3(n5957), .IN4(n5544), .Q(n2576)
         );
  OA22X1 U2943 ( .IN1(n6210), .IN2(n5534), .IN3(n5531), .IN4(n5942), .Q(n2577)
         );
  OAI22X1 U2944 ( .IN1(n5973), .IN2(n5584), .IN3(n5579), .IN4(n2578), .QN(
        N10689) );
  OA22X1 U2945 ( .IN1(n6363), .IN2(n5560), .IN3(n5568), .IN4(n2579), .Q(n2578)
         );
  OA22X1 U2946 ( .IN1(n5551), .IN2(n2580), .IN3(n5958), .IN4(n5544), .Q(n2579)
         );
  OA22X1 U2947 ( .IN1(n6209), .IN2(n5534), .IN3(n5531), .IN4(n5943), .Q(n2580)
         );
  OAI22X1 U2948 ( .IN1(n5974), .IN2(n5584), .IN3(n5579), .IN4(n2581), .QN(
        N10688) );
  OA22X1 U2949 ( .IN1(n6362), .IN2(n5560), .IN3(n5572), .IN4(n2582), .Q(n2581)
         );
  OA22X1 U2950 ( .IN1(n5551), .IN2(n2583), .IN3(n5959), .IN4(n5544), .Q(n2582)
         );
  OA22X1 U2951 ( .IN1(n6208), .IN2(n5534), .IN3(n5531), .IN4(n5944), .Q(n2583)
         );
  OAI22X1 U2952 ( .IN1(n5975), .IN2(n5582), .IN3(n5579), .IN4(n2584), .QN(
        N10687) );
  OA22X1 U2953 ( .IN1(n6308), .IN2(n5560), .IN3(n5571), .IN4(n2585), .Q(n2584)
         );
  OA22X1 U2954 ( .IN1(n5551), .IN2(n2586), .IN3(n5960), .IN4(n5543), .Q(n2585)
         );
  OA22X1 U2955 ( .IN1(n6154), .IN2(n5534), .IN3(n5531), .IN4(n5945), .Q(n2586)
         );
  OAI22X1 U2956 ( .IN1(n5976), .IN2(n5583), .IN3(n5579), .IN4(n2587), .QN(
        N10686) );
  OA22X1 U2957 ( .IN1(n6309), .IN2(n5560), .IN3(n5562), .IN4(n2588), .Q(n2587)
         );
  OA22X1 U2958 ( .IN1(n5551), .IN2(n2589), .IN3(n5961), .IN4(n5543), .Q(n2588)
         );
  OA22X1 U2959 ( .IN1(n6155), .IN2(n5534), .IN3(n5531), .IN4(n5946), .Q(n2589)
         );
  OAI22X1 U2960 ( .IN1(n5977), .IN2(n5584), .IN3(n5579), .IN4(n2590), .QN(
        N10685) );
  OA22X1 U2961 ( .IN1(n6310), .IN2(n5560), .IN3(n5565), .IN4(n2591), .Q(n2590)
         );
  OA22X1 U2962 ( .IN1(n5551), .IN2(n2592), .IN3(n5962), .IN4(n5543), .Q(n2591)
         );
  OA22X1 U2963 ( .IN1(n6156), .IN2(n5535), .IN3(n5531), .IN4(n5947), .Q(n2592)
         );
  OAI22X1 U2964 ( .IN1(n5978), .IN2(n5574), .IN3(n5579), .IN4(n2593), .QN(
        N10684) );
  OA22X1 U2965 ( .IN1(n6311), .IN2(n5560), .IN3(n5572), .IN4(n2594), .Q(n2593)
         );
  OA22X1 U2966 ( .IN1(n5550), .IN2(n2595), .IN3(n5963), .IN4(n5543), .Q(n2594)
         );
  OA22X1 U2967 ( .IN1(n6157), .IN2(n5535), .IN3(n5531), .IN4(n5948), .Q(n2595)
         );
  OAI22X1 U2968 ( .IN1(n5979), .IN2(n5575), .IN3(n5579), .IN4(n2596), .QN(
        N10683) );
  OA22X1 U2969 ( .IN1(n6312), .IN2(n5560), .IN3(n5571), .IN4(n2597), .Q(n2596)
         );
  OA22X1 U2970 ( .IN1(n5550), .IN2(n2598), .IN3(n5964), .IN4(n5543), .Q(n2597)
         );
  OA22X1 U2971 ( .IN1(n6158), .IN2(n5535), .IN3(n5531), .IN4(n5949), .Q(n2598)
         );
  OAI22X1 U2972 ( .IN1(n5980), .IN2(n5573), .IN3(n5579), .IN4(n2599), .QN(
        N10682) );
  OA22X1 U2973 ( .IN1(n6313), .IN2(n5560), .IN3(n5570), .IN4(n2600), .Q(n2599)
         );
  OA22X1 U2974 ( .IN1(n5550), .IN2(n2601), .IN3(n5965), .IN4(n5543), .Q(n2600)
         );
  OA22X1 U2975 ( .IN1(n6159), .IN2(n5535), .IN3(n5531), .IN4(n5950), .Q(n2601)
         );
  OAI22X1 U2976 ( .IN1(n5981), .IN2(n5585), .IN3(n5579), .IN4(n2602), .QN(
        N10681) );
  OA22X1 U2977 ( .IN1(n6314), .IN2(n5560), .IN3(n5571), .IN4(n2603), .Q(n2602)
         );
  OA22X1 U2978 ( .IN1(n5550), .IN2(n2604), .IN3(n5966), .IN4(n5543), .Q(n2603)
         );
  OA22X1 U2979 ( .IN1(n6160), .IN2(n5535), .IN3(n5531), .IN4(n5951), .Q(n2604)
         );
  OAI22X1 U2980 ( .IN1(n6375), .IN2(n5583), .IN3(n5579), .IN4(n2605), .QN(
        N10680) );
  OA22X1 U2981 ( .IN1(n6307), .IN2(n5560), .IN3(n5570), .IN4(n2606), .Q(n2605)
         );
  OA22X1 U2982 ( .IN1(n5550), .IN2(n2607), .IN3(n6221), .IN4(n5543), .Q(n2606)
         );
  OA22X1 U2983 ( .IN1(n6153), .IN2(n5536), .IN3(n5531), .IN4(n6067), .Q(n2607)
         );
  OAI22X1 U2984 ( .IN1(n6372), .IN2(n5583), .IN3(n5579), .IN4(n2608), .QN(
        N10678) );
  OA22X1 U2985 ( .IN1(n6306), .IN2(n5560), .IN3(n5571), .IN4(n2609), .Q(n2608)
         );
  OA22X1 U2986 ( .IN1(n5550), .IN2(n2610), .IN3(n6218), .IN4(n5543), .Q(n2609)
         );
  OA22X1 U2987 ( .IN1(n6152), .IN2(n5536), .IN3(n5531), .IN4(n6064), .Q(n2610)
         );
  OAI22X1 U2988 ( .IN1(n6377), .IN2(n5583), .IN3(n5579), .IN4(n2611), .QN(
        N10676) );
  OA22X1 U2989 ( .IN1(n6422), .IN2(n5560), .IN3(n5572), .IN4(n2612), .Q(n2611)
         );
  OA22X1 U2990 ( .IN1(n5550), .IN2(n2613), .IN3(n6223), .IN4(n5543), .Q(n2612)
         );
  OA22X1 U2991 ( .IN1(n6268), .IN2(n5536), .IN3(n5531), .IN4(n6069), .Q(n2613)
         );
  OAI22X1 U2992 ( .IN1(n6378), .IN2(n5583), .IN3(n5579), .IN4(n2614), .QN(
        N10675) );
  OA22X1 U2993 ( .IN1(n6421), .IN2(n5559), .IN3(n5568), .IN4(n2615), .Q(n2614)
         );
  OA22X1 U2994 ( .IN1(n5550), .IN2(n2616), .IN3(n6224), .IN4(n5543), .Q(n2615)
         );
  OA22X1 U2995 ( .IN1(n6267), .IN2(n5536), .IN3(n5531), .IN4(n6070), .Q(n2616)
         );
  OAI22X1 U2996 ( .IN1(n6379), .IN2(n5583), .IN3(n5579), .IN4(n2617), .QN(
        N10674) );
  OA22X1 U2997 ( .IN1(n6420), .IN2(n5559), .IN3(n5565), .IN4(n2618), .Q(n2617)
         );
  OA22X1 U2998 ( .IN1(n5550), .IN2(n2619), .IN3(n6225), .IN4(n5543), .Q(n2618)
         );
  OA22X1 U2999 ( .IN1(n6266), .IN2(n5536), .IN3(n5531), .IN4(n6071), .Q(n2619)
         );
  OAI22X1 U3000 ( .IN1(n6380), .IN2(n5583), .IN3(n5579), .IN4(n2620), .QN(
        N10673) );
  OA22X1 U3001 ( .IN1(n6419), .IN2(n5559), .IN3(n5570), .IN4(n2621), .Q(n2620)
         );
  OA22X1 U3002 ( .IN1(n5550), .IN2(n2622), .IN3(n6226), .IN4(n5543), .Q(n2621)
         );
  OA22X1 U3003 ( .IN1(n6265), .IN2(n5537), .IN3(n5531), .IN4(n6072), .Q(n2622)
         );
  OAI22X1 U3004 ( .IN1(n6381), .IN2(n5583), .IN3(n5579), .IN4(n2623), .QN(
        N10672) );
  OA22X1 U3005 ( .IN1(n6418), .IN2(n5559), .IN3(n5570), .IN4(n2624), .Q(n2623)
         );
  OA22X1 U3006 ( .IN1(n5550), .IN2(n2625), .IN3(n6227), .IN4(n5543), .Q(n2624)
         );
  OA22X1 U3007 ( .IN1(n6264), .IN2(n5537), .IN3(n5531), .IN4(n6073), .Q(n2625)
         );
  OAI22X1 U3008 ( .IN1(n6382), .IN2(n5582), .IN3(n5579), .IN4(n2626), .QN(
        N10671) );
  OA22X1 U3009 ( .IN1(n6417), .IN2(n5559), .IN3(n5571), .IN4(n2627), .Q(n2626)
         );
  OA22X1 U3010 ( .IN1(n5550), .IN2(n2628), .IN3(n6228), .IN4(n5543), .Q(n2627)
         );
  OA22X1 U3011 ( .IN1(n6263), .IN2(n5537), .IN3(n5531), .IN4(n6074), .Q(n2628)
         );
  OAI22X1 U3012 ( .IN1(n6383), .IN2(n5582), .IN3(n5579), .IN4(n2629), .QN(
        N10670) );
  OA22X1 U3013 ( .IN1(n6416), .IN2(n5559), .IN3(n5572), .IN4(n2630), .Q(n2629)
         );
  OA22X1 U3014 ( .IN1(n5549), .IN2(n2631), .IN3(n6229), .IN4(n5543), .Q(n2630)
         );
  OA22X1 U3015 ( .IN1(n6262), .IN2(n5537), .IN3(n5531), .IN4(n6075), .Q(n2631)
         );
  OAI22X1 U3016 ( .IN1(n6385), .IN2(n5582), .IN3(n5579), .IN4(n2632), .QN(
        N10669) );
  OA22X1 U3017 ( .IN1(n6359), .IN2(n5559), .IN3(n5569), .IN4(n2633), .Q(n2632)
         );
  OA22X1 U3018 ( .IN1(n5549), .IN2(n2634), .IN3(n6231), .IN4(n5543), .Q(n2633)
         );
  OA22X1 U3019 ( .IN1(n6205), .IN2(n5537), .IN3(n5531), .IN4(n6077), .Q(n2634)
         );
  OAI22X1 U3020 ( .IN1(n6386), .IN2(n5582), .IN3(n5579), .IN4(n2635), .QN(
        N10668) );
  OA22X1 U3021 ( .IN1(n6358), .IN2(n5559), .IN3(n5563), .IN4(n2636), .Q(n2635)
         );
  OA22X1 U3022 ( .IN1(n5549), .IN2(n2637), .IN3(n6232), .IN4(n5543), .Q(n2636)
         );
  OA22X1 U3023 ( .IN1(n6204), .IN2(n5538), .IN3(n5531), .IN4(n6078), .Q(n2637)
         );
  OAI22X1 U3024 ( .IN1(n6387), .IN2(n5582), .IN3(n5579), .IN4(n2638), .QN(
        N10667) );
  OA22X1 U3025 ( .IN1(n6357), .IN2(n5559), .IN3(n5565), .IN4(n2639), .Q(n2638)
         );
  OA22X1 U3026 ( .IN1(n5549), .IN2(n2640), .IN3(n6233), .IN4(n5543), .Q(n2639)
         );
  OA22X1 U3027 ( .IN1(n6203), .IN2(n5538), .IN3(n5531), .IN4(n6079), .Q(n2640)
         );
  OAI22X1 U3028 ( .IN1(n6388), .IN2(n5582), .IN3(n5579), .IN4(n2641), .QN(
        N10666) );
  OA22X1 U3029 ( .IN1(n6356), .IN2(n5559), .IN3(n5569), .IN4(n2642), .Q(n2641)
         );
  OA22X1 U3030 ( .IN1(n5549), .IN2(n2643), .IN3(n6234), .IN4(n5543), .Q(n2642)
         );
  OA22X1 U3031 ( .IN1(n6202), .IN2(n5538), .IN3(n5531), .IN4(n6080), .Q(n2643)
         );
  OAI22X1 U3032 ( .IN1(n6389), .IN2(n5582), .IN3(n5579), .IN4(n2644), .QN(
        N10665) );
  OA22X1 U3033 ( .IN1(n6355), .IN2(n5559), .IN3(n5568), .IN4(n2645), .Q(n2644)
         );
  OA22X1 U3034 ( .IN1(n5549), .IN2(n2646), .IN3(n6235), .IN4(n5543), .Q(n2645)
         );
  OA22X1 U3035 ( .IN1(n6201), .IN2(n5538), .IN3(n5530), .IN4(n6081), .Q(n2646)
         );
  OAI22X1 U3036 ( .IN1(n6390), .IN2(n5574), .IN3(n5579), .IN4(n2647), .QN(
        N10664) );
  OA22X1 U3037 ( .IN1(n6354), .IN2(n5559), .IN3(n5566), .IN4(n2648), .Q(n2647)
         );
  OA22X1 U3038 ( .IN1(n5549), .IN2(n2649), .IN3(n6236), .IN4(n5543), .Q(n2648)
         );
  OA22X1 U3039 ( .IN1(n6200), .IN2(n5538), .IN3(n5530), .IN4(n6082), .Q(n2649)
         );
  OAI22X1 U3040 ( .IN1(n6391), .IN2(n5584), .IN3(n5579), .IN4(n2650), .QN(
        N10663) );
  OA22X1 U3041 ( .IN1(n6353), .IN2(n5559), .IN3(n5567), .IN4(n2651), .Q(n2650)
         );
  OA22X1 U3042 ( .IN1(n5549), .IN2(n2652), .IN3(n6237), .IN4(n5543), .Q(n2651)
         );
  OA22X1 U3043 ( .IN1(n6199), .IN2(n5535), .IN3(n5530), .IN4(n6083), .Q(n2652)
         );
  OAI22X1 U3044 ( .IN1(n6400), .IN2(n5575), .IN3(n5579), .IN4(n2653), .QN(
        N10662) );
  OA22X1 U3045 ( .IN1(n6415), .IN2(n5559), .IN3(n5562), .IN4(n2654), .Q(n2653)
         );
  OA22X1 U3046 ( .IN1(n5549), .IN2(n2655), .IN3(n6246), .IN4(n5543), .Q(n2654)
         );
  OA22X1 U3047 ( .IN1(n6261), .IN2(n5536), .IN3(n5530), .IN4(n6092), .Q(n2655)
         );
  OAI22X1 U3048 ( .IN1(n6406), .IN2(n5573), .IN3(n5579), .IN4(n2656), .QN(
        N10661) );
  OA22X1 U3049 ( .IN1(n6414), .IN2(n5558), .IN3(n5563), .IN4(n2657), .Q(n2656)
         );
  OA22X1 U3050 ( .IN1(n5549), .IN2(n2658), .IN3(n6252), .IN4(n5543), .Q(n2657)
         );
  OA22X1 U3051 ( .IN1(n6260), .IN2(n5537), .IN3(n5530), .IN4(n6098), .Q(n2658)
         );
  OAI22X1 U3052 ( .IN1(n6407), .IN2(n5574), .IN3(n5579), .IN4(n2659), .QN(
        N10660) );
  OA22X1 U3053 ( .IN1(n6413), .IN2(n5558), .IN3(n5564), .IN4(n2660), .Q(n2659)
         );
  OA22X1 U3054 ( .IN1(n5549), .IN2(n2661), .IN3(n6253), .IN4(n5543), .Q(n2660)
         );
  OA22X1 U3055 ( .IN1(n6259), .IN2(n5537), .IN3(n5530), .IN4(n6099), .Q(n2661)
         );
  OAI22X1 U3056 ( .IN1(n6408), .IN2(n5585), .IN3(n5579), .IN4(n2662), .QN(
        N10659) );
  OA22X1 U3057 ( .IN1(n6412), .IN2(n5558), .IN3(n5569), .IN4(n2663), .Q(n2662)
         );
  OA22X1 U3058 ( .IN1(n5549), .IN2(n2664), .IN3(n6254), .IN4(n5543), .Q(n2663)
         );
  OA22X1 U3059 ( .IN1(n6258), .IN2(n5532), .IN3(n5530), .IN4(n6100), .Q(n2664)
         );
  OAI22X1 U3060 ( .IN1(n6409), .IN2(n5581), .IN3(n5579), .IN4(n2665), .QN(
        N10658) );
  OA22X1 U3061 ( .IN1(n6411), .IN2(n5558), .IN3(n5563), .IN4(n2666), .Q(n2665)
         );
  OA22X1 U3062 ( .IN1(n5548), .IN2(n2667), .IN3(n6255), .IN4(n5543), .Q(n2666)
         );
  OA22X1 U3063 ( .IN1(n6257), .IN2(n5538), .IN3(n5530), .IN4(n6101), .Q(n2667)
         );
  OAI22X1 U3064 ( .IN1(n6401), .IN2(n5583), .IN3(n5579), .IN4(n2668), .QN(
        N10657) );
  OA22X1 U3065 ( .IN1(n6410), .IN2(n5558), .IN3(n5565), .IN4(n2669), .Q(n2668)
         );
  OA22X1 U3066 ( .IN1(n5548), .IN2(n2670), .IN3(n6247), .IN4(n5543), .Q(n2669)
         );
  OA22X1 U3067 ( .IN1(n6256), .IN2(n5536), .IN3(n5530), .IN4(n6093), .Q(n2670)
         );
  OAI22X1 U3068 ( .IN1(n6399), .IN2(n5582), .IN3(n5579), .IN4(n2671), .QN(
        N10656) );
  OA22X1 U3069 ( .IN1(n6352), .IN2(n5558), .IN3(n5568), .IN4(n2672), .Q(n2671)
         );
  OA22X1 U3070 ( .IN1(n5548), .IN2(n2673), .IN3(n6244), .IN4(n5543), .Q(n2672)
         );
  OA22X1 U3071 ( .IN1(n6198), .IN2(n5534), .IN3(n5530), .IN4(n6090), .Q(n2673)
         );
  OAI22X1 U3072 ( .IN1(n6398), .IN2(n5574), .IN3(n5580), .IN4(n2674), .QN(
        N10655) );
  OA22X1 U3073 ( .IN1(n6402), .IN2(n5558), .IN3(n5562), .IN4(n2675), .Q(n2674)
         );
  OA22X1 U3074 ( .IN1(n5548), .IN2(n2676), .IN3(n6243), .IN4(n5543), .Q(n2675)
         );
  OA22X1 U3075 ( .IN1(n6248), .IN2(n5538), .IN3(n5530), .IN4(n6089), .Q(n2676)
         );
  OAI22X1 U3076 ( .IN1(n6397), .IN2(n5584), .IN3(n5580), .IN4(n2677), .QN(
        N10654) );
  OA22X1 U3077 ( .IN1(n6403), .IN2(n5558), .IN3(n5564), .IN4(n2678), .Q(n2677)
         );
  OA22X1 U3078 ( .IN1(n5548), .IN2(n2679), .IN3(n6242), .IN4(n5543), .Q(n2678)
         );
  OA22X1 U3079 ( .IN1(n6249), .IN2(n5532), .IN3(n5530), .IN4(n6090), .Q(n2679)
         );
  OAI22X1 U3080 ( .IN1(n6396), .IN2(n5573), .IN3(n5580), .IN4(n2680), .QN(
        N10653) );
  OA22X1 U3081 ( .IN1(n6404), .IN2(n5558), .IN3(n5566), .IN4(n2681), .Q(n2680)
         );
  OA22X1 U3082 ( .IN1(n5548), .IN2(n2682), .IN3(n6241), .IN4(n5543), .Q(n2681)
         );
  OA22X1 U3083 ( .IN1(n6250), .IN2(n5538), .IN3(n5530), .IN4(n6088), .Q(n2682)
         );
  OAI22X1 U3084 ( .IN1(n6396), .IN2(n5575), .IN3(n5580), .IN4(n2683), .QN(
        N10652) );
  OA22X1 U3085 ( .IN1(n6405), .IN2(n5558), .IN3(n5563), .IN4(n2684), .Q(n2683)
         );
  OA22X1 U3086 ( .IN1(n5548), .IN2(n2685), .IN3(n6241), .IN4(n5543), .Q(n2684)
         );
  OA22X1 U3087 ( .IN1(n6251), .IN2(n5532), .IN3(n5530), .IN4(n6087), .Q(n2685)
         );
  OAI22X1 U3088 ( .IN1(n6394), .IN2(n5574), .IN3(n5580), .IN4(n2686), .QN(
        N10651) );
  OA22X1 U3089 ( .IN1(n6393), .IN2(n5558), .IN3(n5572), .IN4(n2687), .Q(n2686)
         );
  OA22X1 U3090 ( .IN1(n5548), .IN2(n2688), .IN3(n6240), .IN4(n5543), .Q(n2687)
         );
  OA22X1 U3091 ( .IN1(n6239), .IN2(n5533), .IN3(n5530), .IN4(n6086), .Q(n2688)
         );
  OAI22X1 U3092 ( .IN1(n6361), .IN2(n5585), .IN3(n5580), .IN4(n2689), .QN(
        N10650) );
  OA22X1 U3093 ( .IN1(n6360), .IN2(n5558), .IN3(n5568), .IN4(n2690), .Q(n2689)
         );
  OA22X1 U3094 ( .IN1(n5548), .IN2(n2691), .IN3(n6207), .IN4(n5542), .Q(n2690)
         );
  OA22X1 U3095 ( .IN1(n6206), .IN2(n5534), .IN3(n5530), .IN4(n6053), .Q(n2691)
         );
  OAI22X1 U3096 ( .IN1(n6350), .IN2(n5582), .IN3(n5580), .IN4(n2692), .QN(
        N10649) );
  OA22X1 U3097 ( .IN1(n6351), .IN2(n5558), .IN3(n5568), .IN4(n2693), .Q(n2692)
         );
  OA22X1 U3098 ( .IN1(n5548), .IN2(n2694), .IN3(n6196), .IN4(n5542), .Q(n2693)
         );
  OA22X1 U3099 ( .IN1(n6197), .IN2(n5535), .IN3(n5530), .IN4(n6042), .Q(n2694)
         );
  OAI22X1 U3100 ( .IN1(n6395), .IN2(n5583), .IN3(n5580), .IN4(n2695), .QN(
        N10648) );
  OA22X1 U3101 ( .IN1(n6392), .IN2(n5558), .IN3(n5569), .IN4(n2696), .Q(n2695)
         );
  OA22X1 U3102 ( .IN1(n5548), .IN2(n2697), .IN3(n6241), .IN4(n5542), .Q(n2696)
         );
  OA22X1 U3103 ( .IN1(n6238), .IN2(n5537), .IN3(n5530), .IN4(n6088), .Q(n2697)
         );
  OAI22X1 U3104 ( .IN1(n6423), .IN2(n5581), .IN3(n5580), .IN4(n2698), .QN(
        N10647) );
  OA22X1 U3105 ( .IN1(n6423), .IN2(n5557), .IN3(n5570), .IN4(n2699), .Q(n2698)
         );
  OA22X1 U3106 ( .IN1(n5548), .IN2(n2700), .IN3(n6269), .IN4(n5542), .Q(n2699)
         );
  OA22X1 U3107 ( .IN1(n6269), .IN2(n5532), .IN3(n5530), .IN4(n6115), .Q(n2700)
         );
  OAI22X1 U3108 ( .IN1(n6424), .IN2(n5574), .IN3(n5580), .IN4(n2701), .QN(
        N10646) );
  OA22X1 U3109 ( .IN1(n6424), .IN2(n5557), .IN3(n5565), .IN4(n2702), .Q(n2701)
         );
  OA22X1 U3110 ( .IN1(n5547), .IN2(n2703), .IN3(n6270), .IN4(n5542), .Q(n2702)
         );
  OA22X1 U3111 ( .IN1(n6270), .IN2(n5533), .IN3(n5530), .IN4(n6116), .Q(n2703)
         );
  OAI22X1 U3112 ( .IN1(n6425), .IN2(n5584), .IN3(n5580), .IN4(n2704), .QN(
        N10645) );
  OA22X1 U3113 ( .IN1(n6425), .IN2(n5557), .IN3(n5570), .IN4(n2705), .Q(n2704)
         );
  OA22X1 U3114 ( .IN1(n5547), .IN2(n2706), .IN3(n6271), .IN4(n5542), .Q(n2705)
         );
  OA22X1 U3115 ( .IN1(n6271), .IN2(n5534), .IN3(n5530), .IN4(n6117), .Q(n2706)
         );
  OAI22X1 U3116 ( .IN1(n6426), .IN2(n5575), .IN3(n5580), .IN4(n2707), .QN(
        N10644) );
  OA22X1 U3117 ( .IN1(n6426), .IN2(n5557), .IN3(n5565), .IN4(n2708), .Q(n2707)
         );
  OA22X1 U3118 ( .IN1(n5547), .IN2(n2709), .IN3(n6272), .IN4(n5542), .Q(n2708)
         );
  OA22X1 U3119 ( .IN1(n6272), .IN2(n5535), .IN3(n5530), .IN4(n6118), .Q(n2709)
         );
  OAI22X1 U3120 ( .IN1(n6427), .IN2(n5581), .IN3(n5580), .IN4(n2710), .QN(
        N10643) );
  OA22X1 U3121 ( .IN1(n6427), .IN2(n5557), .IN3(n5571), .IN4(n2711), .Q(n2710)
         );
  OA22X1 U3122 ( .IN1(n5547), .IN2(n2712), .IN3(n6273), .IN4(n5542), .Q(n2711)
         );
  OA22X1 U3123 ( .IN1(n6273), .IN2(n5538), .IN3(n5530), .IN4(n6119), .Q(n2712)
         );
  OAI22X1 U3124 ( .IN1(n6428), .IN2(n5581), .IN3(n5580), .IN4(n2713), .QN(
        N10642) );
  OA22X1 U3125 ( .IN1(n6428), .IN2(n5557), .IN3(n5570), .IN4(n2714), .Q(n2713)
         );
  OA22X1 U3126 ( .IN1(n5547), .IN2(n2715), .IN3(n6274), .IN4(n5542), .Q(n2714)
         );
  OA22X1 U3127 ( .IN1(n6274), .IN2(n5538), .IN3(n5530), .IN4(n6120), .Q(n2715)
         );
  OAI22X1 U3128 ( .IN1(n6429), .IN2(n5581), .IN3(n5580), .IN4(n2716), .QN(
        N10641) );
  OA22X1 U3129 ( .IN1(n6429), .IN2(n5557), .IN3(n5572), .IN4(n2717), .Q(n2716)
         );
  OA22X1 U3130 ( .IN1(n5547), .IN2(n2718), .IN3(n6275), .IN4(n5542), .Q(n2717)
         );
  OA22X1 U3131 ( .IN1(n6275), .IN2(n5532), .IN3(n5530), .IN4(n6121), .Q(n2718)
         );
  OAI22X1 U3132 ( .IN1(n6430), .IN2(n5581), .IN3(n5580), .IN4(n2719), .QN(
        N10640) );
  OA22X1 U3133 ( .IN1(n6430), .IN2(n5557), .IN3(n5567), .IN4(n2720), .Q(n2719)
         );
  OA22X1 U3134 ( .IN1(n5547), .IN2(n2721), .IN3(n6276), .IN4(n5542), .Q(n2720)
         );
  OA22X1 U3135 ( .IN1(n6276), .IN2(n5533), .IN3(n5530), .IN4(n6122), .Q(n2721)
         );
  OAI22X1 U3136 ( .IN1(n6431), .IN2(n5581), .IN3(n5580), .IN4(n2722), .QN(
        N10639) );
  OA22X1 U3137 ( .IN1(n6431), .IN2(n5557), .IN3(n5567), .IN4(n2723), .Q(n2722)
         );
  OA22X1 U3138 ( .IN1(n5547), .IN2(n2724), .IN3(n6277), .IN4(n5542), .Q(n2723)
         );
  OA22X1 U3139 ( .IN1(n6277), .IN2(n5534), .IN3(n5530), .IN4(n6123), .Q(n2724)
         );
  OAI22X1 U3140 ( .IN1(n6432), .IN2(n5581), .IN3(n5580), .IN4(n2725), .QN(
        N10638) );
  OA22X1 U3141 ( .IN1(n6432), .IN2(n5557), .IN3(n5564), .IN4(n2726), .Q(n2725)
         );
  OA22X1 U3142 ( .IN1(n5547), .IN2(n2727), .IN3(n6278), .IN4(n5542), .Q(n2726)
         );
  OA22X1 U3143 ( .IN1(n6278), .IN2(n5534), .IN3(n5530), .IN4(n6124), .Q(n2727)
         );
  OAI22X1 U3144 ( .IN1(n6433), .IN2(n5581), .IN3(n5580), .IN4(n2728), .QN(
        N10637) );
  OA22X1 U3145 ( .IN1(n6433), .IN2(n5557), .IN3(n5566), .IN4(n2729), .Q(n2728)
         );
  OA22X1 U3146 ( .IN1(n5547), .IN2(n2730), .IN3(n6279), .IN4(n5542), .Q(n2729)
         );
  OA22X1 U3147 ( .IN1(n6279), .IN2(n5532), .IN3(n5530), .IN4(n6125), .Q(n2730)
         );
  OAI22X1 U3148 ( .IN1(n6434), .IN2(n5581), .IN3(n5580), .IN4(n2731), .QN(
        N10636) );
  OA22X1 U3149 ( .IN1(n6434), .IN2(n5557), .IN3(n5562), .IN4(n2732), .Q(n2731)
         );
  OA22X1 U3150 ( .IN1(n5547), .IN2(n2733), .IN3(n6280), .IN4(n5542), .Q(n2732)
         );
  OA22X1 U3151 ( .IN1(n6280), .IN2(n5533), .IN3(n5530), .IN4(n6126), .Q(n2733)
         );
  OAI22X1 U3152 ( .IN1(n6435), .IN2(n5583), .IN3(n5580), .IN4(n2734), .QN(
        N10635) );
  OA22X1 U3153 ( .IN1(n6435), .IN2(n5557), .IN3(n5563), .IN4(n2735), .Q(n2734)
         );
  OA22X1 U3154 ( .IN1(n5547), .IN2(n2736), .IN3(n6281), .IN4(n5542), .Q(n2735)
         );
  OA22X1 U3155 ( .IN1(n6281), .IN2(n5534), .IN3(n5530), .IN4(n6127), .Q(n2736)
         );
  OAI22X1 U3156 ( .IN1(n6436), .IN2(n5581), .IN3(n5580), .IN4(n2737), .QN(
        N10634) );
  OA22X1 U3157 ( .IN1(n6436), .IN2(n5557), .IN3(n5562), .IN4(n2738), .Q(n2737)
         );
  OA22X1 U3158 ( .IN1(n5546), .IN2(n2739), .IN3(n6282), .IN4(n5542), .Q(n2738)
         );
  OA22X1 U3159 ( .IN1(n6282), .IN2(n5538), .IN3(n5530), .IN4(n6128), .Q(n2739)
         );
  OAI22X1 U3160 ( .IN1(n6437), .IN2(n5584), .IN3(n5580), .IN4(n2740), .QN(
        N10633) );
  OA22X1 U3161 ( .IN1(n6437), .IN2(n5556), .IN3(n5562), .IN4(n2741), .Q(n2740)
         );
  OA22X1 U3162 ( .IN1(n5546), .IN2(n2742), .IN3(n6283), .IN4(n5542), .Q(n2741)
         );
  OA22X1 U3163 ( .IN1(n6283), .IN2(n5537), .IN3(n5530), .IN4(n6129), .Q(n2742)
         );
  OAI22X1 U3164 ( .IN1(n6438), .IN2(n5575), .IN3(n5580), .IN4(n2743), .QN(
        N10632) );
  OA22X1 U3165 ( .IN1(n6438), .IN2(n5556), .IN3(n5562), .IN4(n2744), .Q(n2743)
         );
  OA22X1 U3166 ( .IN1(n5546), .IN2(n2745), .IN3(n6284), .IN4(n5542), .Q(n2744)
         );
  OA22X1 U3167 ( .IN1(n6284), .IN2(n5533), .IN3(n5530), .IN4(n6130), .Q(n2745)
         );
  OAI22X1 U3168 ( .IN1(n6439), .IN2(n5582), .IN3(n5580), .IN4(n2746), .QN(
        N10631) );
  OA22X1 U3169 ( .IN1(n6439), .IN2(n5556), .IN3(n5562), .IN4(n2747), .Q(n2746)
         );
  OA22X1 U3170 ( .IN1(n5546), .IN2(n2748), .IN3(n6285), .IN4(n5542), .Q(n2747)
         );
  OA22X1 U3171 ( .IN1(n6285), .IN2(n5532), .IN3(n5530), .IN4(n6131), .Q(n2748)
         );
  OAI22X1 U3172 ( .IN1(n6440), .IN2(n5573), .IN3(n5580), .IN4(n2749), .QN(
        N10630) );
  OA22X1 U3173 ( .IN1(n6440), .IN2(n5556), .IN3(n5562), .IN4(n2750), .Q(n2749)
         );
  OA22X1 U3174 ( .IN1(n5546), .IN2(n2751), .IN3(n6286), .IN4(n5542), .Q(n2750)
         );
  OA22X1 U3175 ( .IN1(n6286), .IN2(n5535), .IN3(n5530), .IN4(n6132), .Q(n2751)
         );
  OAI22X1 U3176 ( .IN1(n6441), .IN2(n5573), .IN3(n5580), .IN4(n2752), .QN(
        N10629) );
  OA22X1 U3177 ( .IN1(n6441), .IN2(n5556), .IN3(n5563), .IN4(n2753), .Q(n2752)
         );
  OA22X1 U3178 ( .IN1(n5546), .IN2(n2754), .IN3(n6287), .IN4(n5542), .Q(n2753)
         );
  OA22X1 U3179 ( .IN1(n6287), .IN2(n5533), .IN3(n5530), .IN4(n6133), .Q(n2754)
         );
  OAI22X1 U3180 ( .IN1(n6442), .IN2(n5573), .IN3(n5580), .IN4(n2755), .QN(
        N10628) );
  OA22X1 U3181 ( .IN1(n6442), .IN2(n5556), .IN3(n5563), .IN4(n2756), .Q(n2755)
         );
  OA22X1 U3182 ( .IN1(n5546), .IN2(n2757), .IN3(n6288), .IN4(n5542), .Q(n2756)
         );
  OA22X1 U3183 ( .IN1(n6288), .IN2(n5533), .IN3(n5275), .IN4(n6134), .Q(n2757)
         );
  OAI22X1 U3184 ( .IN1(n6443), .IN2(n5582), .IN3(n5580), .IN4(n2758), .QN(
        N10626) );
  OA22X1 U3185 ( .IN1(n6443), .IN2(n5556), .IN3(n5563), .IN4(n2759), .Q(n2758)
         );
  OA22X1 U3186 ( .IN1(n5546), .IN2(n2760), .IN3(n6289), .IN4(n5542), .Q(n2759)
         );
  OA22X1 U3187 ( .IN1(n6289), .IN2(n5534), .IN3(n5275), .IN4(n6135), .Q(n2760)
         );
  OAI22X1 U3188 ( .IN1(n6444), .IN2(n5585), .IN3(n5580), .IN4(n2761), .QN(
        N10625) );
  OA22X1 U3189 ( .IN1(n6444), .IN2(n5556), .IN3(n5563), .IN4(n2762), .Q(n2761)
         );
  OA22X1 U3190 ( .IN1(n5546), .IN2(n2763), .IN3(n6290), .IN4(n5542), .Q(n2762)
         );
  OA22X1 U3191 ( .IN1(n6290), .IN2(n5535), .IN3(n5275), .IN4(n6136), .Q(n2763)
         );
  OAI22X1 U3192 ( .IN1(n6445), .IN2(n5584), .IN3(n5580), .IN4(n2764), .QN(
        N10624) );
  OA22X1 U3193 ( .IN1(n6445), .IN2(n5556), .IN3(n5563), .IN4(n2765), .Q(n2764)
         );
  OA22X1 U3194 ( .IN1(n5546), .IN2(n2766), .IN3(n6291), .IN4(n5542), .Q(n2765)
         );
  OA22X1 U3195 ( .IN1(n6291), .IN2(n5536), .IN3(n5275), .IN4(n6137), .Q(n2766)
         );
  OAI22X1 U3196 ( .IN1(n6446), .IN2(n5573), .IN3(n5580), .IN4(n2767), .QN(
        N10623) );
  OA22X1 U3197 ( .IN1(n6446), .IN2(n5556), .IN3(n5564), .IN4(n2768), .Q(n2767)
         );
  OA22X1 U3198 ( .IN1(n5546), .IN2(n2769), .IN3(n6292), .IN4(n5542), .Q(n2768)
         );
  OA22X1 U3199 ( .IN1(n6292), .IN2(n5536), .IN3(n5275), .IN4(n6138), .Q(n2769)
         );
  OAI22X1 U3200 ( .IN1(n6447), .IN2(n5575), .IN3(n5580), .IN4(n2770), .QN(
        N10622) );
  OA22X1 U3201 ( .IN1(n6447), .IN2(n5556), .IN3(n5564), .IN4(n2771), .Q(n2770)
         );
  OA22X1 U3202 ( .IN1(n5546), .IN2(n2772), .IN3(n6293), .IN4(n5542), .Q(n2771)
         );
  OA22X1 U3203 ( .IN1(n6293), .IN2(n5535), .IN3(n5275), .IN4(n6139), .Q(n2772)
         );
  OAI22X1 U3204 ( .IN1(n6448), .IN2(n5581), .IN3(n5580), .IN4(n2773), .QN(
        N10621) );
  OA22X1 U3205 ( .IN1(n6448), .IN2(n5556), .IN3(n5564), .IN4(n2774), .Q(n2773)
         );
  OA22X1 U3206 ( .IN1(n5545), .IN2(n2775), .IN3(n6294), .IN4(n5542), .Q(n2774)
         );
  OA22X1 U3207 ( .IN1(n6294), .IN2(n5534), .IN3(n5275), .IN4(n6140), .Q(n2775)
         );
  OAI22X1 U3208 ( .IN1(n6449), .IN2(n5581), .IN3(n5580), .IN4(n2776), .QN(
        N10620) );
  OA22X1 U3209 ( .IN1(n6449), .IN2(n5556), .IN3(n5564), .IN4(n2777), .Q(n2776)
         );
  OA22X1 U3210 ( .IN1(n5545), .IN2(n2778), .IN3(n6295), .IN4(n5542), .Q(n2777)
         );
  OA22X1 U3211 ( .IN1(n6295), .IN2(n5537), .IN3(n5275), .IN4(n6141), .Q(n2778)
         );
  OAI22X1 U3212 ( .IN1(n6450), .IN2(n5573), .IN3(n5580), .IN4(n2779), .QN(
        N10619) );
  OA22X1 U3213 ( .IN1(n6450), .IN2(n5556), .IN3(n5564), .IN4(n2780), .Q(n2779)
         );
  OA22X1 U3214 ( .IN1(n5545), .IN2(n2781), .IN3(n6296), .IN4(n5542), .Q(n2780)
         );
  OA22X1 U3215 ( .IN1(n6296), .IN2(n5538), .IN3(n5275), .IN4(n6142), .Q(n2781)
         );
  OAI22X1 U3216 ( .IN1(n6451), .IN2(n5573), .IN3(n5580), .IN4(n2782), .QN(
        N10618) );
  OA22X1 U3217 ( .IN1(n6451), .IN2(n5555), .IN3(n5565), .IN4(n2783), .Q(n2782)
         );
  OA22X1 U3218 ( .IN1(n5545), .IN2(n2784), .IN3(n6297), .IN4(n5542), .Q(n2783)
         );
  OA22X1 U3219 ( .IN1(n6297), .IN2(n5536), .IN3(n5275), .IN4(n6143), .Q(n2784)
         );
  OAI22X1 U3220 ( .IN1(n6452), .IN2(n5583), .IN3(n5580), .IN4(n2785), .QN(
        N10617) );
  OA22X1 U3221 ( .IN1(n6452), .IN2(n5555), .IN3(n5565), .IN4(n2786), .Q(n2785)
         );
  OA22X1 U3222 ( .IN1(n5545), .IN2(n2787), .IN3(n6298), .IN4(n5542), .Q(n2786)
         );
  OA22X1 U3223 ( .IN1(n6298), .IN2(n5536), .IN3(n5275), .IN4(n6144), .Q(n2787)
         );
  OAI22X1 U3224 ( .IN1(n6453), .IN2(n5582), .IN3(n5580), .IN4(n2788), .QN(
        N10616) );
  OA22X1 U3225 ( .IN1(n6453), .IN2(n5555), .IN3(n5565), .IN4(n2789), .Q(n2788)
         );
  OA22X1 U3226 ( .IN1(n5545), .IN2(n2790), .IN3(n6299), .IN4(n5542), .Q(n2789)
         );
  OA22X1 U3227 ( .IN1(n6299), .IN2(n5537), .IN3(n5275), .IN4(n6145), .Q(n2790)
         );
  OAI22X1 U3228 ( .IN1(n6454), .IN2(n5575), .IN3(n5577), .IN4(n2791), .QN(
        N10615) );
  OA22X1 U3229 ( .IN1(n6454), .IN2(n5555), .IN3(n5565), .IN4(n2792), .Q(n2791)
         );
  OA22X1 U3230 ( .IN1(n5545), .IN2(n2793), .IN3(n6300), .IN4(n5542), .Q(n2792)
         );
  OA22X1 U3231 ( .IN1(n6300), .IN2(n5535), .IN3(n5275), .IN4(n6146), .Q(n2793)
         );
  OA22X1 U3233 ( .IN1(n6320), .IN2(n5555), .IN3(n5565), .IN4(n2795), .Q(n2794)
         );
  OA22X1 U3237 ( .IN1(n6321), .IN2(n5555), .IN3(n5566), .IN4(n2798), .Q(n2797)
         );
  OA22X1 U3241 ( .IN1(n6322), .IN2(n5555), .IN3(n5566), .IN4(n2801), .Q(n2800)
         );
  OA22X1 U3245 ( .IN1(n6323), .IN2(n5555), .IN3(n5566), .IN4(n2804), .Q(n2803)
         );
  OA22X1 U3249 ( .IN1(n6324), .IN2(n5555), .IN3(n5566), .IN4(n2807), .Q(n2806)
         );
  OA22X1 U3253 ( .IN1(n6325), .IN2(n5555), .IN3(n5566), .IN4(n2810), .Q(n2809)
         );
  OA22X1 U3257 ( .IN1(n6326), .IN2(n5555), .IN3(n5567), .IN4(n2813), .Q(n2812)
         );
  OA22X1 U3261 ( .IN1(n6327), .IN2(n5555), .IN3(n5567), .IN4(n2816), .Q(n2815)
         );
  OA22X1 U3265 ( .IN1(n6328), .IN2(n5555), .IN3(n5567), .IN4(n2819), .Q(n2818)
         );
  OA22X1 U3269 ( .IN1(n6329), .IN2(n5555), .IN3(n5567), .IN4(n2822), .Q(n2821)
         );
  OA22X1 U3273 ( .IN1(n6330), .IN2(n5554), .IN3(n5567), .IN4(n2825), .Q(n2824)
         );
  OA22X1 U3277 ( .IN1(n6331), .IN2(n5554), .IN3(n5568), .IN4(n2828), .Q(n2827)
         );
  OA22X1 U3281 ( .IN1(n6332), .IN2(n5554), .IN3(n5568), .IN4(n2831), .Q(n2830)
         );
  OA22X1 U3285 ( .IN1(n6333), .IN2(n5554), .IN3(n5568), .IN4(n2834), .Q(n2833)
         );
  OA22X1 U3289 ( .IN1(n6334), .IN2(n5554), .IN3(n5568), .IN4(n2837), .Q(n2836)
         );
  OA22X1 U3293 ( .IN1(n6335), .IN2(n5554), .IN3(n5568), .IN4(n2840), .Q(n2839)
         );
  OA22X1 U3297 ( .IN1(n6336), .IN2(n5554), .IN3(n5569), .IN4(n2843), .Q(n2842)
         );
  OA22X1 U3301 ( .IN1(n6337), .IN2(n5554), .IN3(n5569), .IN4(n2846), .Q(n2845)
         );
  OA22X1 U3305 ( .IN1(n6338), .IN2(n5554), .IN3(n5569), .IN4(n2849), .Q(n2848)
         );
  OA22X1 U3309 ( .IN1(n6339), .IN2(n5554), .IN3(n5569), .IN4(n2852), .Q(n2851)
         );
  OA22X1 U3313 ( .IN1(n6340), .IN2(n5554), .IN3(n5569), .IN4(n2855), .Q(n2854)
         );
  OA22X1 U3317 ( .IN1(n6341), .IN2(n5554), .IN3(n5565), .IN4(n2858), .Q(n2857)
         );
  OA22X1 U3321 ( .IN1(n6342), .IN2(n5554), .IN3(n5570), .IN4(n2861), .Q(n2860)
         );
  OA22X1 U3325 ( .IN1(n6343), .IN2(n5554), .IN3(n5571), .IN4(n2864), .Q(n2863)
         );
  OA22X1 U3329 ( .IN1(n6344), .IN2(n5553), .IN3(n5567), .IN4(n2867), .Q(n2866)
         );
  OA22X1 U3333 ( .IN1(n6345), .IN2(n5553), .IN3(n5564), .IN4(n2870), .Q(n2869)
         );
  OA22X1 U3337 ( .IN1(n6346), .IN2(n5553), .IN3(n5566), .IN4(n2873), .Q(n2872)
         );
  OA22X1 U3341 ( .IN1(n6315), .IN2(n5553), .IN3(n5567), .IN4(n2876), .Q(n2875)
         );
  OA22X1 U3345 ( .IN1(n6316), .IN2(n5553), .IN3(n5562), .IN4(n2879), .Q(n2878)
         );
  OA22X1 U3349 ( .IN1(n6317), .IN2(n5553), .IN3(n5563), .IN4(n2882), .Q(n2881)
         );
  OA22X1 U3353 ( .IN1(n6318), .IN2(n5553), .IN3(n5564), .IN4(n2885), .Q(n2884)
         );
  OA22X1 U3357 ( .IN1(n6319), .IN2(n5553), .IN3(n5569), .IN4(n2888), .Q(n2887)
         );
  OAI22X1 U3360 ( .IN1(n6455), .IN2(n5573), .IN3(n5576), .IN4(n2890), .QN(
        N10582) );
  OA22X1 U3361 ( .IN1(n6455), .IN2(n5553), .IN3(n5568), .IN4(n2891), .Q(n2890)
         );
  OA22X1 U3362 ( .IN1(n5545), .IN2(n2892), .IN3(n6301), .IN4(n5541), .Q(n2891)
         );
  OA22X1 U3363 ( .IN1(n6301), .IN2(n5537), .IN3(n5275), .IN4(n6147), .Q(n2892)
         );
  OAI22X1 U3364 ( .IN1(n6456), .IN2(n5585), .IN3(n5577), .IN4(n2893), .QN(
        N10581) );
  OA22X1 U3365 ( .IN1(n6456), .IN2(n5553), .IN3(n5566), .IN4(n2894), .Q(n2893)
         );
  OA22X1 U3366 ( .IN1(n5545), .IN2(n2895), .IN3(n6302), .IN4(n5541), .Q(n2894)
         );
  OA22X1 U3367 ( .IN1(n6302), .IN2(n5536), .IN3(n5275), .IN4(n6148), .Q(n2895)
         );
  OAI22X1 U3368 ( .IN1(n6457), .IN2(n5583), .IN3(n5576), .IN4(n2896), .QN(
        N10580) );
  OA22X1 U3369 ( .IN1(n6457), .IN2(n5553), .IN3(n5566), .IN4(n2897), .Q(n2896)
         );
  OA22X1 U3370 ( .IN1(n5545), .IN2(n2898), .IN3(n6303), .IN4(n5541), .Q(n2897)
         );
  OA22X1 U3371 ( .IN1(n6303), .IN2(n5538), .IN3(n5275), .IN4(n6149), .Q(n2898)
         );
  OAI22X1 U3372 ( .IN1(n6458), .IN2(n5574), .IN3(n5577), .IN4(n2899), .QN(
        N10579) );
  OA22X1 U3373 ( .IN1(n6458), .IN2(n5553), .IN3(n5570), .IN4(n2900), .Q(n2899)
         );
  OA22X1 U3374 ( .IN1(n5545), .IN2(n2901), .IN3(n6304), .IN4(n5541), .Q(n2900)
         );
  OA22X1 U3375 ( .IN1(n6304), .IN2(n5532), .IN3(n5275), .IN4(n6150), .Q(n2901)
         );
  OAI22X1 U3376 ( .IN1(n6459), .IN2(n5573), .IN3(n5576), .IN4(n2902), .QN(
        N10578) );
  OA22X1 U3377 ( .IN1(n6459), .IN2(n5553), .IN3(n5570), .IN4(n2903), .Q(n2902)
         );
  OA22X1 U3378 ( .IN1(n5545), .IN2(n2904), .IN3(n6305), .IN4(n5541), .Q(n2903)
         );
  OA22X1 U3379 ( .IN1(n6305), .IN2(n5533), .IN3(n5530), .IN4(n6151), .Q(n2904)
         );
  NAND4X0 U3380 ( .IN1(n2905), .IN2(n5553), .IN3(n2906), .IN4(n5541), .QN(
        decodedVector_o[7]) );
  NAND4X0 U3382 ( .IN1(decodedPacketValid[4]), .IN2(N2173), .IN3(N2172), .IN4(
        n2908), .QN(n2529) );
  NAND4X0 U3383 ( .IN1(decodedPacketValid[7]), .IN2(N8581), .IN3(N8580), .IN4(
        n2909), .QN(n2523) );
  NAND4X0 U3384 ( .IN1(decodedPacketValid[6]), .IN2(N6445), .IN3(N6444), .IN4(
        n2910), .QN(n2525) );
  NAND4X0 U3385 ( .IN1(decodedPacketValid[3]), .IN2(N1069), .IN3(N1068), .IN4(
        N1070), .QN(n2905) );
  OA22X1 U3403 ( .IN1(n5856), .IN2(n5503), .IN3(n5507), .IN4(n2929), .Q(n2928)
         );
  OAI22X1 U3406 ( .IN1(n6384), .IN2(n5527), .IN3(n5519), .IN4(n2931), .QN(
        N10571) );
  OA22X1 U3407 ( .IN1(n6349), .IN2(n5503), .IN3(n5513), .IN4(n2932), .Q(n2931)
         );
  OA22X1 U3408 ( .IN1(n5494), .IN2(n2933), .IN3(n6230), .IN4(n5486), .Q(n2932)
         );
  OA22X1 U3409 ( .IN1(n6195), .IN2(n5473), .IN3(n5273), .IN4(n6076), .Q(n2933)
         );
  OAI22X1 U3410 ( .IN1(n6376), .IN2(n5527), .IN3(n5519), .IN4(n2934), .QN(
        N10570) );
  OA22X1 U3411 ( .IN1(n6348), .IN2(n5503), .IN3(n5507), .IN4(n2935), .Q(n2934)
         );
  OA22X1 U3412 ( .IN1(n5494), .IN2(n2936), .IN3(n6222), .IN4(n5486), .Q(n2935)
         );
  OA22X1 U3413 ( .IN1(n6194), .IN2(n5473), .IN3(n5472), .IN4(n6068), .Q(n2936)
         );
  OAI22X1 U3414 ( .IN1(n6372), .IN2(n5527), .IN3(n5519), .IN4(n2937), .QN(
        N10569) );
  OA22X1 U3415 ( .IN1(n6374), .IN2(n5503), .IN3(n5504), .IN4(n2938), .Q(n2937)
         );
  OA22X1 U3416 ( .IN1(n5494), .IN2(n2939), .IN3(n6218), .IN4(n5486), .Q(n2938)
         );
  OA22X1 U3417 ( .IN1(n6220), .IN2(n5473), .IN3(n5472), .IN4(n6065), .Q(n2939)
         );
  OA22X1 U3419 ( .IN1(n6371), .IN2(n5503), .IN3(n5511), .IN4(n2941), .Q(n2940)
         );
  OAI22X1 U3422 ( .IN1(n6373), .IN2(n5527), .IN3(n5519), .IN4(n2943), .QN(
        N10567) );
  OA22X1 U3423 ( .IN1(n6370), .IN2(n5503), .IN3(n5510), .IN4(n2944), .Q(n2943)
         );
  OA22X1 U3424 ( .IN1(n5494), .IN2(n2945), .IN3(n6219), .IN4(n5486), .Q(n2944)
         );
  OA22X1 U3425 ( .IN1(n6216), .IN2(n5473), .IN3(n5472), .IN4(n6065), .Q(n2945)
         );
  OAI22X1 U3426 ( .IN1(n6396), .IN2(n5527), .IN3(n5520), .IN4(n2946), .QN(
        N10566) );
  OA22X1 U3427 ( .IN1(n6347), .IN2(n5503), .IN3(n5509), .IN4(n2947), .Q(n2946)
         );
  OA22X1 U3428 ( .IN1(n5493), .IN2(n2948), .IN3(n6245), .IN4(n5486), .Q(n2947)
         );
  OA22X1 U3429 ( .IN1(n6193), .IN2(n5473), .IN3(n5472), .IN4(n6091), .Q(n2948)
         );
  OAI22X1 U3430 ( .IN1(n5967), .IN2(n5527), .IN3(n5520), .IN4(n2949), .QN(
        N10565) );
  OA22X1 U3431 ( .IN1(n6369), .IN2(n5503), .IN3(n5504), .IN4(n2950), .Q(n2949)
         );
  OA22X1 U3432 ( .IN1(n5493), .IN2(n2951), .IN3(n5952), .IN4(n5486), .Q(n2950)
         );
  OA22X1 U3433 ( .IN1(n6215), .IN2(n5474), .IN3(n5472), .IN4(n5937), .Q(n2951)
         );
  OAI22X1 U3434 ( .IN1(n5968), .IN2(n5526), .IN3(n5520), .IN4(n2952), .QN(
        N10564) );
  OA22X1 U3435 ( .IN1(n6368), .IN2(n5503), .IN3(n5505), .IN4(n2953), .Q(n2952)
         );
  OA22X1 U3436 ( .IN1(n5493), .IN2(n2954), .IN3(n5953), .IN4(n5486), .Q(n2953)
         );
  OA22X1 U3437 ( .IN1(n6214), .IN2(n5474), .IN3(n5472), .IN4(n5938), .Q(n2954)
         );
  OAI22X1 U3438 ( .IN1(n5969), .IN2(n5526), .IN3(n5520), .IN4(n2955), .QN(
        N10563) );
  OA22X1 U3439 ( .IN1(n6367), .IN2(n5503), .IN3(n5506), .IN4(n2956), .Q(n2955)
         );
  OA22X1 U3440 ( .IN1(n5493), .IN2(n2957), .IN3(n5954), .IN4(n5486), .Q(n2956)
         );
  OA22X1 U3441 ( .IN1(n6213), .IN2(n5474), .IN3(n5472), .IN4(n5939), .Q(n2957)
         );
  OAI22X1 U3442 ( .IN1(n5970), .IN2(n5526), .IN3(n5520), .IN4(n2958), .QN(
        N10562) );
  OA22X1 U3443 ( .IN1(n6366), .IN2(n5503), .IN3(n5514), .IN4(n2959), .Q(n2958)
         );
  OA22X1 U3444 ( .IN1(n5493), .IN2(n2960), .IN3(n5955), .IN4(n5486), .Q(n2959)
         );
  OA22X1 U3445 ( .IN1(n6212), .IN2(n5474), .IN3(n5472), .IN4(n5940), .Q(n2960)
         );
  OAI22X1 U3446 ( .IN1(n5971), .IN2(n5526), .IN3(n5520), .IN4(n2961), .QN(
        N10561) );
  OA22X1 U3447 ( .IN1(n6365), .IN2(n5502), .IN3(n5508), .IN4(n2962), .Q(n2961)
         );
  OA22X1 U3448 ( .IN1(n5493), .IN2(n2963), .IN3(n5956), .IN4(n5486), .Q(n2962)
         );
  OA22X1 U3449 ( .IN1(n6211), .IN2(n5474), .IN3(n5472), .IN4(n5941), .Q(n2963)
         );
  OAI22X1 U3450 ( .IN1(n5972), .IN2(n5526), .IN3(n5520), .IN4(n2964), .QN(
        N10560) );
  OA22X1 U3451 ( .IN1(n6364), .IN2(n5502), .IN3(n5511), .IN4(n2965), .Q(n2964)
         );
  OA22X1 U3452 ( .IN1(n5493), .IN2(n2966), .IN3(n5957), .IN4(n5486), .Q(n2965)
         );
  OA22X1 U3453 ( .IN1(n6210), .IN2(n5475), .IN3(n5472), .IN4(n5942), .Q(n2966)
         );
  OAI22X1 U3454 ( .IN1(n5973), .IN2(n5526), .IN3(n5520), .IN4(n2967), .QN(
        N10559) );
  OA22X1 U3455 ( .IN1(n6363), .IN2(n5502), .IN3(n5510), .IN4(n2968), .Q(n2967)
         );
  OA22X1 U3456 ( .IN1(n5493), .IN2(n2969), .IN3(n5958), .IN4(n5486), .Q(n2968)
         );
  OA22X1 U3457 ( .IN1(n6209), .IN2(n5475), .IN3(n5472), .IN4(n5943), .Q(n2969)
         );
  OAI22X1 U3458 ( .IN1(n5974), .IN2(n5526), .IN3(n5520), .IN4(n2970), .QN(
        N10558) );
  OA22X1 U3459 ( .IN1(n6362), .IN2(n5502), .IN3(n5514), .IN4(n2971), .Q(n2970)
         );
  OA22X1 U3460 ( .IN1(n5493), .IN2(n2972), .IN3(n5959), .IN4(n5486), .Q(n2971)
         );
  OA22X1 U3461 ( .IN1(n6208), .IN2(n5475), .IN3(n5472), .IN4(n5944), .Q(n2972)
         );
  OAI22X1 U3462 ( .IN1(n5975), .IN2(n5525), .IN3(n5520), .IN4(n2973), .QN(
        N10557) );
  OA22X1 U3463 ( .IN1(n6308), .IN2(n5502), .IN3(n5513), .IN4(n2974), .Q(n2973)
         );
  OA22X1 U3464 ( .IN1(n5493), .IN2(n2975), .IN3(n5960), .IN4(n5485), .Q(n2974)
         );
  OA22X1 U3465 ( .IN1(n6154), .IN2(n5475), .IN3(n5472), .IN4(n5945), .Q(n2975)
         );
  OAI22X1 U3466 ( .IN1(n5976), .IN2(n5525), .IN3(n5520), .IN4(n2976), .QN(
        N10556) );
  OA22X1 U3467 ( .IN1(n6309), .IN2(n5502), .IN3(n5504), .IN4(n2977), .Q(n2976)
         );
  OA22X1 U3468 ( .IN1(n5493), .IN2(n2978), .IN3(n5961), .IN4(n5485), .Q(n2977)
         );
  OA22X1 U3469 ( .IN1(n6155), .IN2(n5475), .IN3(n5472), .IN4(n5946), .Q(n2978)
         );
  OAI22X1 U3470 ( .IN1(n5977), .IN2(n5525), .IN3(n5520), .IN4(n2979), .QN(
        N10555) );
  OA22X1 U3471 ( .IN1(n6310), .IN2(n5502), .IN3(n5507), .IN4(n2980), .Q(n2979)
         );
  OA22X1 U3472 ( .IN1(n5493), .IN2(n2981), .IN3(n5962), .IN4(n5485), .Q(n2980)
         );
  OA22X1 U3473 ( .IN1(n6156), .IN2(n5476), .IN3(n5472), .IN4(n5947), .Q(n2981)
         );
  OAI22X1 U3474 ( .IN1(n5978), .IN2(n5525), .IN3(n5520), .IN4(n2982), .QN(
        N10554) );
  OA22X1 U3475 ( .IN1(n6311), .IN2(n5502), .IN3(n5514), .IN4(n2983), .Q(n2982)
         );
  OA22X1 U3476 ( .IN1(n5492), .IN2(n2984), .IN3(n5963), .IN4(n5485), .Q(n2983)
         );
  OA22X1 U3477 ( .IN1(n6157), .IN2(n5476), .IN3(n5472), .IN4(n5948), .Q(n2984)
         );
  OAI22X1 U3478 ( .IN1(n5979), .IN2(n5525), .IN3(n5520), .IN4(n2985), .QN(
        N10553) );
  OA22X1 U3479 ( .IN1(n6312), .IN2(n5502), .IN3(n5513), .IN4(n2986), .Q(n2985)
         );
  OA22X1 U3480 ( .IN1(n5492), .IN2(n2987), .IN3(n5964), .IN4(n5485), .Q(n2986)
         );
  OA22X1 U3481 ( .IN1(n6158), .IN2(n5476), .IN3(n5472), .IN4(n5949), .Q(n2987)
         );
  OAI22X1 U3482 ( .IN1(n5980), .IN2(n5525), .IN3(n5520), .IN4(n2988), .QN(
        N10552) );
  OA22X1 U3483 ( .IN1(n6313), .IN2(n5502), .IN3(n5512), .IN4(n2989), .Q(n2988)
         );
  OA22X1 U3484 ( .IN1(n5492), .IN2(n2990), .IN3(n5965), .IN4(n5485), .Q(n2989)
         );
  OA22X1 U3485 ( .IN1(n6159), .IN2(n5476), .IN3(n5472), .IN4(n5950), .Q(n2990)
         );
  OAI22X1 U3486 ( .IN1(n5981), .IN2(n5525), .IN3(n5520), .IN4(n2991), .QN(
        N10551) );
  OA22X1 U3487 ( .IN1(n6314), .IN2(n5502), .IN3(n5513), .IN4(n2992), .Q(n2991)
         );
  OA22X1 U3488 ( .IN1(n5492), .IN2(n2993), .IN3(n5966), .IN4(n5485), .Q(n2992)
         );
  OA22X1 U3489 ( .IN1(n6160), .IN2(n5476), .IN3(n5472), .IN4(n5951), .Q(n2993)
         );
  OAI22X1 U3490 ( .IN1(n6375), .IN2(n5524), .IN3(n5520), .IN4(n2994), .QN(
        N10550) );
  OA22X1 U3491 ( .IN1(n6307), .IN2(n5502), .IN3(n5512), .IN4(n2995), .Q(n2994)
         );
  OA22X1 U3492 ( .IN1(n5492), .IN2(n2996), .IN3(n6221), .IN4(n5485), .Q(n2995)
         );
  OA22X1 U3493 ( .IN1(n6153), .IN2(n5477), .IN3(n5472), .IN4(n6067), .Q(n2996)
         );
  OAI22X1 U3494 ( .IN1(n6372), .IN2(n5524), .IN3(n5520), .IN4(n2997), .QN(
        N10548) );
  OA22X1 U3495 ( .IN1(n6306), .IN2(n5502), .IN3(n5513), .IN4(n2998), .Q(n2997)
         );
  OA22X1 U3496 ( .IN1(n5492), .IN2(n2999), .IN3(n6218), .IN4(n5485), .Q(n2998)
         );
  OA22X1 U3497 ( .IN1(n6152), .IN2(n5477), .IN3(n5472), .IN4(n6064), .Q(n2999)
         );
  OAI22X1 U3498 ( .IN1(n6377), .IN2(n5524), .IN3(n5520), .IN4(n3000), .QN(
        N10546) );
  OA22X1 U3499 ( .IN1(n6422), .IN2(n5502), .IN3(n5514), .IN4(n3001), .Q(n3000)
         );
  OA22X1 U3500 ( .IN1(n5492), .IN2(n3002), .IN3(n6223), .IN4(n5485), .Q(n3001)
         );
  OA22X1 U3501 ( .IN1(n6268), .IN2(n5477), .IN3(n5472), .IN4(n6069), .Q(n3002)
         );
  OAI22X1 U3502 ( .IN1(n6378), .IN2(n5524), .IN3(n5520), .IN4(n3003), .QN(
        N10545) );
  OA22X1 U3503 ( .IN1(n6421), .IN2(n5501), .IN3(n5510), .IN4(n3004), .Q(n3003)
         );
  OA22X1 U3504 ( .IN1(n5492), .IN2(n3005), .IN3(n6224), .IN4(n5485), .Q(n3004)
         );
  OA22X1 U3505 ( .IN1(n6267), .IN2(n5477), .IN3(n5472), .IN4(n6070), .Q(n3005)
         );
  OAI22X1 U3506 ( .IN1(n6379), .IN2(n5524), .IN3(n5520), .IN4(n3006), .QN(
        N10544) );
  OA22X1 U3507 ( .IN1(n6420), .IN2(n5501), .IN3(n5507), .IN4(n3007), .Q(n3006)
         );
  OA22X1 U3508 ( .IN1(n5492), .IN2(n3008), .IN3(n6225), .IN4(n5485), .Q(n3007)
         );
  OA22X1 U3509 ( .IN1(n6266), .IN2(n5477), .IN3(n5472), .IN4(n6071), .Q(n3008)
         );
  OAI22X1 U3510 ( .IN1(n6380), .IN2(n5524), .IN3(n5520), .IN4(n3009), .QN(
        N10543) );
  OA22X1 U3511 ( .IN1(n6419), .IN2(n5501), .IN3(n5512), .IN4(n3010), .Q(n3009)
         );
  OA22X1 U3512 ( .IN1(n5492), .IN2(n3011), .IN3(n6226), .IN4(n5485), .Q(n3010)
         );
  OA22X1 U3513 ( .IN1(n6265), .IN2(n5478), .IN3(n5472), .IN4(n6072), .Q(n3011)
         );
  OAI22X1 U3514 ( .IN1(n6381), .IN2(n5524), .IN3(n5520), .IN4(n3012), .QN(
        N10542) );
  OA22X1 U3515 ( .IN1(n6418), .IN2(n5501), .IN3(n5512), .IN4(n3013), .Q(n3012)
         );
  OA22X1 U3516 ( .IN1(n5492), .IN2(n3014), .IN3(n6227), .IN4(n5485), .Q(n3013)
         );
  OA22X1 U3517 ( .IN1(n6264), .IN2(n5478), .IN3(n5472), .IN4(n6073), .Q(n3014)
         );
  OAI22X1 U3518 ( .IN1(n6382), .IN2(n5523), .IN3(n5520), .IN4(n3015), .QN(
        N10541) );
  OA22X1 U3519 ( .IN1(n6417), .IN2(n5501), .IN3(n5513), .IN4(n3016), .Q(n3015)
         );
  OA22X1 U3520 ( .IN1(n5492), .IN2(n3017), .IN3(n6228), .IN4(n5485), .Q(n3016)
         );
  OA22X1 U3521 ( .IN1(n6263), .IN2(n5478), .IN3(n5472), .IN4(n6074), .Q(n3017)
         );
  OAI22X1 U3522 ( .IN1(n6383), .IN2(n5523), .IN3(n5520), .IN4(n3018), .QN(
        N10540) );
  OA22X1 U3523 ( .IN1(n6416), .IN2(n5501), .IN3(n5514), .IN4(n3019), .Q(n3018)
         );
  OA22X1 U3524 ( .IN1(n5491), .IN2(n3020), .IN3(n6229), .IN4(n5485), .Q(n3019)
         );
  OA22X1 U3525 ( .IN1(n6262), .IN2(n5478), .IN3(n5472), .IN4(n6075), .Q(n3020)
         );
  OAI22X1 U3526 ( .IN1(n6385), .IN2(n5523), .IN3(n5520), .IN4(n3021), .QN(
        N10539) );
  OA22X1 U3527 ( .IN1(n6359), .IN2(n5501), .IN3(n5511), .IN4(n3022), .Q(n3021)
         );
  OA22X1 U3528 ( .IN1(n5491), .IN2(n3023), .IN3(n6231), .IN4(n5485), .Q(n3022)
         );
  OA22X1 U3529 ( .IN1(n6205), .IN2(n5478), .IN3(n5472), .IN4(n6077), .Q(n3023)
         );
  OAI22X1 U3530 ( .IN1(n6386), .IN2(n5523), .IN3(n5520), .IN4(n3024), .QN(
        N10538) );
  OA22X1 U3531 ( .IN1(n6358), .IN2(n5501), .IN3(n5505), .IN4(n3025), .Q(n3024)
         );
  OA22X1 U3532 ( .IN1(n5491), .IN2(n3026), .IN3(n6232), .IN4(n5485), .Q(n3025)
         );
  OA22X1 U3533 ( .IN1(n6204), .IN2(n5479), .IN3(n5472), .IN4(n6078), .Q(n3026)
         );
  OAI22X1 U3534 ( .IN1(n6387), .IN2(n5523), .IN3(n5520), .IN4(n3027), .QN(
        N10537) );
  OA22X1 U3535 ( .IN1(n6357), .IN2(n5501), .IN3(n5507), .IN4(n3028), .Q(n3027)
         );
  OA22X1 U3536 ( .IN1(n5491), .IN2(n3029), .IN3(n6233), .IN4(n5485), .Q(n3028)
         );
  OA22X1 U3537 ( .IN1(n6203), .IN2(n5479), .IN3(n5472), .IN4(n6079), .Q(n3029)
         );
  OAI22X1 U3538 ( .IN1(n6388), .IN2(n5523), .IN3(n5520), .IN4(n3030), .QN(
        N10536) );
  OA22X1 U3539 ( .IN1(n6356), .IN2(n5501), .IN3(n5511), .IN4(n3031), .Q(n3030)
         );
  OA22X1 U3540 ( .IN1(n5491), .IN2(n3032), .IN3(n6234), .IN4(n5485), .Q(n3031)
         );
  OA22X1 U3541 ( .IN1(n6202), .IN2(n5479), .IN3(n5472), .IN4(n6080), .Q(n3032)
         );
  OAI22X1 U3542 ( .IN1(n6389), .IN2(n5523), .IN3(n5520), .IN4(n3033), .QN(
        N10535) );
  OA22X1 U3543 ( .IN1(n6355), .IN2(n5501), .IN3(n5510), .IN4(n3034), .Q(n3033)
         );
  OA22X1 U3544 ( .IN1(n5491), .IN2(n3035), .IN3(n6235), .IN4(n5485), .Q(n3034)
         );
  OA22X1 U3545 ( .IN1(n6201), .IN2(n5479), .IN3(n5471), .IN4(n6081), .Q(n3035)
         );
  OAI22X1 U3546 ( .IN1(n6390), .IN2(n5522), .IN3(n5520), .IN4(n3036), .QN(
        N10534) );
  OA22X1 U3547 ( .IN1(n6354), .IN2(n5501), .IN3(n5508), .IN4(n3037), .Q(n3036)
         );
  OA22X1 U3548 ( .IN1(n5491), .IN2(n3038), .IN3(n6236), .IN4(n5485), .Q(n3037)
         );
  OA22X1 U3549 ( .IN1(n6200), .IN2(n5479), .IN3(n5471), .IN4(n6082), .Q(n3038)
         );
  OAI22X1 U3550 ( .IN1(n6391), .IN2(n5522), .IN3(n5520), .IN4(n3039), .QN(
        N10533) );
  OA22X1 U3551 ( .IN1(n6353), .IN2(n5501), .IN3(n5509), .IN4(n3040), .Q(n3039)
         );
  OA22X1 U3552 ( .IN1(n5491), .IN2(n3041), .IN3(n6237), .IN4(n5485), .Q(n3040)
         );
  OA22X1 U3553 ( .IN1(n6199), .IN2(n5480), .IN3(n5471), .IN4(n6083), .Q(n3041)
         );
  OAI22X1 U3554 ( .IN1(n6400), .IN2(n5522), .IN3(n5520), .IN4(n3042), .QN(
        N10532) );
  OA22X1 U3555 ( .IN1(n6415), .IN2(n5501), .IN3(n5504), .IN4(n3043), .Q(n3042)
         );
  OA22X1 U3556 ( .IN1(n5491), .IN2(n3044), .IN3(n6246), .IN4(n5485), .Q(n3043)
         );
  OA22X1 U3557 ( .IN1(n6261), .IN2(n5475), .IN3(n5471), .IN4(n6092), .Q(n3044)
         );
  OAI22X1 U3558 ( .IN1(n6406), .IN2(n5522), .IN3(n5520), .IN4(n3045), .QN(
        N10531) );
  OA22X1 U3559 ( .IN1(n6414), .IN2(n5500), .IN3(n5505), .IN4(n3046), .Q(n3045)
         );
  OA22X1 U3560 ( .IN1(n5491), .IN2(n3047), .IN3(n6252), .IN4(n5485), .Q(n3046)
         );
  OA22X1 U3561 ( .IN1(n6260), .IN2(n5478), .IN3(n5471), .IN4(n6098), .Q(n3047)
         );
  OAI22X1 U3562 ( .IN1(n6407), .IN2(n5522), .IN3(n5520), .IN4(n3048), .QN(
        N10530) );
  OA22X1 U3563 ( .IN1(n6413), .IN2(n5500), .IN3(n5506), .IN4(n3049), .Q(n3048)
         );
  OA22X1 U3564 ( .IN1(n5491), .IN2(n3050), .IN3(n6253), .IN4(n5485), .Q(n3049)
         );
  OA22X1 U3565 ( .IN1(n6259), .IN2(n5476), .IN3(n5471), .IN4(n6099), .Q(n3050)
         );
  OAI22X1 U3566 ( .IN1(n6408), .IN2(n5522), .IN3(n5520), .IN4(n3051), .QN(
        N10529) );
  OA22X1 U3567 ( .IN1(n6412), .IN2(n5500), .IN3(n5511), .IN4(n3052), .Q(n3051)
         );
  OA22X1 U3568 ( .IN1(n5491), .IN2(n3053), .IN3(n6254), .IN4(n5485), .Q(n3052)
         );
  OA22X1 U3569 ( .IN1(n6258), .IN2(n5473), .IN3(n5471), .IN4(n6100), .Q(n3053)
         );
  OAI22X1 U3570 ( .IN1(n6409), .IN2(n5522), .IN3(n5520), .IN4(n3054), .QN(
        N10528) );
  OA22X1 U3571 ( .IN1(n6411), .IN2(n5500), .IN3(n5505), .IN4(n3055), .Q(n3054)
         );
  OA22X1 U3572 ( .IN1(n5490), .IN2(n3056), .IN3(n6255), .IN4(n5485), .Q(n3055)
         );
  OA22X1 U3573 ( .IN1(n6257), .IN2(n5480), .IN3(n5471), .IN4(n6101), .Q(n3056)
         );
  OAI22X1 U3574 ( .IN1(n6401), .IN2(n5522), .IN3(n5520), .IN4(n3057), .QN(
        N10527) );
  OA22X1 U3575 ( .IN1(n6410), .IN2(n5500), .IN3(n5507), .IN4(n3058), .Q(n3057)
         );
  OA22X1 U3576 ( .IN1(n5490), .IN2(n3059), .IN3(n6247), .IN4(n5485), .Q(n3058)
         );
  OA22X1 U3577 ( .IN1(n6256), .IN2(n5480), .IN3(n5471), .IN4(n6093), .Q(n3059)
         );
  OAI22X1 U3578 ( .IN1(n6399), .IN2(n5515), .IN3(n5520), .IN4(n3060), .QN(
        N10526) );
  OA22X1 U3579 ( .IN1(n6352), .IN2(n5500), .IN3(n5510), .IN4(n3061), .Q(n3060)
         );
  OA22X1 U3580 ( .IN1(n5490), .IN2(n3062), .IN3(n6244), .IN4(n5485), .Q(n3061)
         );
  OA22X1 U3581 ( .IN1(n6198), .IN2(n5480), .IN3(n5471), .IN4(n6090), .Q(n3062)
         );
  OAI22X1 U3582 ( .IN1(n6398), .IN2(n5516), .IN3(n5521), .IN4(n3063), .QN(
        N10525) );
  OA22X1 U3583 ( .IN1(n6402), .IN2(n5500), .IN3(n5504), .IN4(n3064), .Q(n3063)
         );
  OA22X1 U3584 ( .IN1(n5490), .IN2(n3065), .IN3(n6243), .IN4(n5485), .Q(n3064)
         );
  OA22X1 U3585 ( .IN1(n6248), .IN2(n5480), .IN3(n5471), .IN4(n6089), .Q(n3065)
         );
  OAI22X1 U3586 ( .IN1(n6397), .IN2(n5523), .IN3(n5521), .IN4(n3066), .QN(
        N10524) );
  OA22X1 U3587 ( .IN1(n6403), .IN2(n5500), .IN3(n5506), .IN4(n3067), .Q(n3066)
         );
  OA22X1 U3588 ( .IN1(n5490), .IN2(n3068), .IN3(n6242), .IN4(n5485), .Q(n3067)
         );
  OA22X1 U3589 ( .IN1(n6249), .IN2(n5480), .IN3(n5471), .IN4(n6089), .Q(n3068)
         );
  OAI22X1 U3590 ( .IN1(n6396), .IN2(n5523), .IN3(n5521), .IN4(n3069), .QN(
        N10523) );
  OA22X1 U3591 ( .IN1(n6404), .IN2(n5500), .IN3(n5508), .IN4(n3070), .Q(n3069)
         );
  OA22X1 U3592 ( .IN1(n5490), .IN2(n3071), .IN3(n6241), .IN4(n5485), .Q(n3070)
         );
  OA22X1 U3593 ( .IN1(n6250), .IN2(n5480), .IN3(n5471), .IN4(n6088), .Q(n3071)
         );
  OAI22X1 U3594 ( .IN1(n6397), .IN2(n5524), .IN3(n5521), .IN4(n3072), .QN(
        N10522) );
  OA22X1 U3595 ( .IN1(n6405), .IN2(n5500), .IN3(n5505), .IN4(n3073), .Q(n3072)
         );
  OA22X1 U3596 ( .IN1(n5490), .IN2(n3074), .IN3(n6244), .IN4(n5485), .Q(n3073)
         );
  OA22X1 U3597 ( .IN1(n6251), .IN2(n5478), .IN3(n5471), .IN4(n6087), .Q(n3074)
         );
  OAI22X1 U3598 ( .IN1(n6394), .IN2(n5515), .IN3(n5521), .IN4(n3075), .QN(
        N10521) );
  OA22X1 U3599 ( .IN1(n6393), .IN2(n5500), .IN3(n5514), .IN4(n3076), .Q(n3075)
         );
  OA22X1 U3600 ( .IN1(n5490), .IN2(n3077), .IN3(n6240), .IN4(n5485), .Q(n3076)
         );
  OA22X1 U3601 ( .IN1(n6239), .IN2(n5474), .IN3(n5471), .IN4(n6086), .Q(n3077)
         );
  OAI22X1 U3602 ( .IN1(n6361), .IN2(n5516), .IN3(n5521), .IN4(n3078), .QN(
        N10520) );
  OA22X1 U3603 ( .IN1(n6360), .IN2(n5500), .IN3(n5510), .IN4(n3079), .Q(n3078)
         );
  OA22X1 U3604 ( .IN1(n5490), .IN2(n3080), .IN3(n6207), .IN4(n5484), .Q(n3079)
         );
  OA22X1 U3605 ( .IN1(n6206), .IN2(n5475), .IN3(n5471), .IN4(n6053), .Q(n3080)
         );
  OAI22X1 U3606 ( .IN1(n6350), .IN2(n5527), .IN3(n5521), .IN4(n3081), .QN(
        N10519) );
  OA22X1 U3607 ( .IN1(n6351), .IN2(n5500), .IN3(n5510), .IN4(n3082), .Q(n3081)
         );
  OA22X1 U3608 ( .IN1(n5490), .IN2(n3083), .IN3(n6196), .IN4(n5484), .Q(n3082)
         );
  OA22X1 U3609 ( .IN1(n6197), .IN2(n5476), .IN3(n5471), .IN4(n6042), .Q(n3083)
         );
  OAI22X1 U3610 ( .IN1(n6395), .IN2(n5522), .IN3(n5521), .IN4(n3084), .QN(
        N10518) );
  OA22X1 U3611 ( .IN1(n6392), .IN2(n5500), .IN3(n5511), .IN4(n3085), .Q(n3084)
         );
  OA22X1 U3612 ( .IN1(n5490), .IN2(n3086), .IN3(n6242), .IN4(n5484), .Q(n3085)
         );
  OA22X1 U3613 ( .IN1(n6238), .IN2(n5476), .IN3(n5471), .IN4(n6087), .Q(n3086)
         );
  OAI22X1 U3614 ( .IN1(n6423), .IN2(n5523), .IN3(n5521), .IN4(n3087), .QN(
        N10517) );
  OA22X1 U3615 ( .IN1(n6423), .IN2(n5499), .IN3(n5512), .IN4(n3088), .Q(n3087)
         );
  OA22X1 U3616 ( .IN1(n5490), .IN2(n3089), .IN3(n6269), .IN4(n5484), .Q(n3088)
         );
  OA22X1 U3617 ( .IN1(n6269), .IN2(n5478), .IN3(n5471), .IN4(n6115), .Q(n3089)
         );
  OAI22X1 U3618 ( .IN1(n6424), .IN2(n5524), .IN3(n5521), .IN4(n3090), .QN(
        N10516) );
  OA22X1 U3619 ( .IN1(n6424), .IN2(n5499), .IN3(n5507), .IN4(n3091), .Q(n3090)
         );
  OA22X1 U3620 ( .IN1(n5489), .IN2(n3092), .IN3(n6270), .IN4(n5484), .Q(n3091)
         );
  OA22X1 U3621 ( .IN1(n6270), .IN2(n5475), .IN3(n5471), .IN4(n6116), .Q(n3092)
         );
  OAI22X1 U3622 ( .IN1(n6425), .IN2(n5525), .IN3(n5521), .IN4(n3093), .QN(
        N10515) );
  OA22X1 U3623 ( .IN1(n6425), .IN2(n5499), .IN3(n5512), .IN4(n3094), .Q(n3093)
         );
  OA22X1 U3624 ( .IN1(n5489), .IN2(n3095), .IN3(n6271), .IN4(n5484), .Q(n3094)
         );
  OA22X1 U3625 ( .IN1(n6271), .IN2(n5477), .IN3(n5471), .IN4(n6117), .Q(n3095)
         );
  OAI22X1 U3626 ( .IN1(n6426), .IN2(n5526), .IN3(n5521), .IN4(n3096), .QN(
        N10514) );
  OA22X1 U3627 ( .IN1(n6426), .IN2(n5499), .IN3(n5507), .IN4(n3097), .Q(n3096)
         );
  OA22X1 U3628 ( .IN1(n5489), .IN2(n3098), .IN3(n6272), .IN4(n5484), .Q(n3097)
         );
  OA22X1 U3629 ( .IN1(n6272), .IN2(n5473), .IN3(n5471), .IN4(n6118), .Q(n3098)
         );
  OAI22X1 U3630 ( .IN1(n6427), .IN2(n5525), .IN3(n5521), .IN4(n3099), .QN(
        N10513) );
  OA22X1 U3631 ( .IN1(n6427), .IN2(n5499), .IN3(n5513), .IN4(n3100), .Q(n3099)
         );
  OA22X1 U3632 ( .IN1(n5489), .IN2(n3101), .IN3(n6273), .IN4(n5484), .Q(n3100)
         );
  OA22X1 U3633 ( .IN1(n6273), .IN2(n5477), .IN3(n5471), .IN4(n6119), .Q(n3101)
         );
  OAI22X1 U3634 ( .IN1(n6428), .IN2(n5526), .IN3(n5521), .IN4(n3102), .QN(
        N10512) );
  OA22X1 U3635 ( .IN1(n6428), .IN2(n5499), .IN3(n5512), .IN4(n3103), .Q(n3102)
         );
  OA22X1 U3636 ( .IN1(n5489), .IN2(n3104), .IN3(n6274), .IN4(n5484), .Q(n3103)
         );
  OA22X1 U3637 ( .IN1(n6274), .IN2(n5473), .IN3(n5471), .IN4(n6120), .Q(n3104)
         );
  OAI22X1 U3638 ( .IN1(n6429), .IN2(n5527), .IN3(n5521), .IN4(n3105), .QN(
        N10511) );
  OA22X1 U3639 ( .IN1(n6429), .IN2(n5499), .IN3(n5514), .IN4(n3106), .Q(n3105)
         );
  OA22X1 U3640 ( .IN1(n5489), .IN2(n3107), .IN3(n6275), .IN4(n5484), .Q(n3106)
         );
  OA22X1 U3641 ( .IN1(n6275), .IN2(n5479), .IN3(n5471), .IN4(n6121), .Q(n3107)
         );
  OAI22X1 U3642 ( .IN1(n6430), .IN2(n5522), .IN3(n5521), .IN4(n3108), .QN(
        N10510) );
  OA22X1 U3643 ( .IN1(n6430), .IN2(n5499), .IN3(n5509), .IN4(n3109), .Q(n3108)
         );
  OA22X1 U3644 ( .IN1(n5489), .IN2(n3110), .IN3(n6276), .IN4(n5484), .Q(n3109)
         );
  OA22X1 U3645 ( .IN1(n6276), .IN2(n5480), .IN3(n5471), .IN4(n6122), .Q(n3110)
         );
  OAI22X1 U3646 ( .IN1(n6431), .IN2(n5524), .IN3(n5521), .IN4(n3111), .QN(
        N10509) );
  OA22X1 U3647 ( .IN1(n6431), .IN2(n5499), .IN3(n5509), .IN4(n3112), .Q(n3111)
         );
  OA22X1 U3648 ( .IN1(n5489), .IN2(n3113), .IN3(n6277), .IN4(n5484), .Q(n3112)
         );
  OA22X1 U3649 ( .IN1(n6277), .IN2(n5480), .IN3(n5471), .IN4(n6123), .Q(n3113)
         );
  OAI22X1 U3650 ( .IN1(n6432), .IN2(n5525), .IN3(n5521), .IN4(n3114), .QN(
        N10508) );
  OA22X1 U3651 ( .IN1(n6432), .IN2(n5499), .IN3(n5506), .IN4(n3115), .Q(n3114)
         );
  OA22X1 U3652 ( .IN1(n5489), .IN2(n3116), .IN3(n6278), .IN4(n5484), .Q(n3115)
         );
  OA22X1 U3653 ( .IN1(n6278), .IN2(n5479), .IN3(n5471), .IN4(n6124), .Q(n3116)
         );
  OAI22X1 U3654 ( .IN1(n6433), .IN2(n5526), .IN3(n5521), .IN4(n3117), .QN(
        N10507) );
  OA22X1 U3655 ( .IN1(n6433), .IN2(n5499), .IN3(n5508), .IN4(n3118), .Q(n3117)
         );
  OA22X1 U3656 ( .IN1(n5489), .IN2(n3119), .IN3(n6279), .IN4(n5484), .Q(n3118)
         );
  OA22X1 U3657 ( .IN1(n6279), .IN2(n5479), .IN3(n5471), .IN4(n6125), .Q(n3119)
         );
  OAI22X1 U3658 ( .IN1(n6434), .IN2(n5523), .IN3(n5521), .IN4(n3120), .QN(
        N10506) );
  OA22X1 U3659 ( .IN1(n6434), .IN2(n5499), .IN3(n5504), .IN4(n3121), .Q(n3120)
         );
  OA22X1 U3660 ( .IN1(n5489), .IN2(n3122), .IN3(n6280), .IN4(n5484), .Q(n3121)
         );
  OA22X1 U3661 ( .IN1(n6280), .IN2(n5480), .IN3(n5471), .IN4(n6126), .Q(n3122)
         );
  OAI22X1 U3662 ( .IN1(n6435), .IN2(n5527), .IN3(n5521), .IN4(n3123), .QN(
        N10505) );
  OA22X1 U3663 ( .IN1(n6435), .IN2(n5499), .IN3(n5505), .IN4(n3124), .Q(n3123)
         );
  OA22X1 U3664 ( .IN1(n5489), .IN2(n3125), .IN3(n6281), .IN4(n5484), .Q(n3124)
         );
  OA22X1 U3665 ( .IN1(n6281), .IN2(n5477), .IN3(n5471), .IN4(n6127), .Q(n3125)
         );
  OAI22X1 U3666 ( .IN1(n6436), .IN2(n5516), .IN3(n5521), .IN4(n3126), .QN(
        N10504) );
  OA22X1 U3667 ( .IN1(n6436), .IN2(n5499), .IN3(n5504), .IN4(n3127), .Q(n3126)
         );
  OA22X1 U3668 ( .IN1(n5488), .IN2(n3128), .IN3(n6282), .IN4(n5484), .Q(n3127)
         );
  OA22X1 U3669 ( .IN1(n6282), .IN2(n5474), .IN3(n5471), .IN4(n6128), .Q(n3128)
         );
  OAI22X1 U3670 ( .IN1(n6437), .IN2(n5524), .IN3(n5521), .IN4(n3129), .QN(
        N10503) );
  OA22X1 U3671 ( .IN1(n6437), .IN2(n5498), .IN3(n5504), .IN4(n3130), .Q(n3129)
         );
  OA22X1 U3672 ( .IN1(n5488), .IN2(n3131), .IN3(n6283), .IN4(n5484), .Q(n3130)
         );
  OA22X1 U3673 ( .IN1(n6283), .IN2(n5474), .IN3(n5471), .IN4(n6129), .Q(n3131)
         );
  OAI22X1 U3674 ( .IN1(n6438), .IN2(n5515), .IN3(n5521), .IN4(n3132), .QN(
        N10502) );
  OA22X1 U3675 ( .IN1(n6438), .IN2(n5498), .IN3(n5504), .IN4(n3133), .Q(n3132)
         );
  OA22X1 U3676 ( .IN1(n5488), .IN2(n3134), .IN3(n6284), .IN4(n5484), .Q(n3133)
         );
  OA22X1 U3677 ( .IN1(n6284), .IN2(n5477), .IN3(n5471), .IN4(n6130), .Q(n3134)
         );
  OAI22X1 U3678 ( .IN1(n6439), .IN2(n5522), .IN3(n5521), .IN4(n3135), .QN(
        N10501) );
  OA22X1 U3679 ( .IN1(n6439), .IN2(n5498), .IN3(n5504), .IN4(n3136), .Q(n3135)
         );
  OA22X1 U3680 ( .IN1(n5488), .IN2(n3137), .IN3(n6285), .IN4(n5484), .Q(n3136)
         );
  OA22X1 U3681 ( .IN1(n6285), .IN2(n5473), .IN3(n5471), .IN4(n6131), .Q(n3137)
         );
  OAI22X1 U3682 ( .IN1(n6440), .IN2(n5523), .IN3(n5521), .IN4(n3138), .QN(
        N10500) );
  OA22X1 U3683 ( .IN1(n6440), .IN2(n5498), .IN3(n5504), .IN4(n3139), .Q(n3138)
         );
  OA22X1 U3684 ( .IN1(n5488), .IN2(n3140), .IN3(n6286), .IN4(n5484), .Q(n3139)
         );
  OA22X1 U3685 ( .IN1(n6286), .IN2(n5476), .IN3(n5471), .IN4(n6132), .Q(n3140)
         );
  OAI22X1 U3686 ( .IN1(n6441), .IN2(n5522), .IN3(n5521), .IN4(n3141), .QN(
        N10499) );
  OA22X1 U3687 ( .IN1(n6441), .IN2(n5498), .IN3(n5505), .IN4(n3142), .Q(n3141)
         );
  OA22X1 U3688 ( .IN1(n5488), .IN2(n3143), .IN3(n6287), .IN4(n5484), .Q(n3142)
         );
  OA22X1 U3689 ( .IN1(n6287), .IN2(n5475), .IN3(n5471), .IN4(n6133), .Q(n3143)
         );
  OAI22X1 U3690 ( .IN1(n6442), .IN2(n5523), .IN3(n5521), .IN4(n3144), .QN(
        N10498) );
  OA22X1 U3691 ( .IN1(n6442), .IN2(n5498), .IN3(n5505), .IN4(n3145), .Q(n3144)
         );
  OA22X1 U3692 ( .IN1(n5488), .IN2(n3146), .IN3(n6288), .IN4(n5484), .Q(n3145)
         );
  OA22X1 U3693 ( .IN1(n6288), .IN2(n5473), .IN3(n5273), .IN4(n6134), .Q(n3146)
         );
  OAI22X1 U3694 ( .IN1(n6443), .IN2(n5524), .IN3(n5521), .IN4(n3147), .QN(
        N10496) );
  OA22X1 U3695 ( .IN1(n6443), .IN2(n5498), .IN3(n5505), .IN4(n3148), .Q(n3147)
         );
  OA22X1 U3696 ( .IN1(n5488), .IN2(n3149), .IN3(n6289), .IN4(n5484), .Q(n3148)
         );
  OA22X1 U3697 ( .IN1(n6289), .IN2(n5479), .IN3(n5273), .IN4(n6135), .Q(n3149)
         );
  OAI22X1 U3698 ( .IN1(n6444), .IN2(n5525), .IN3(n5521), .IN4(n3150), .QN(
        N10495) );
  OA22X1 U3699 ( .IN1(n6444), .IN2(n5498), .IN3(n5505), .IN4(n3151), .Q(n3150)
         );
  OA22X1 U3700 ( .IN1(n5488), .IN2(n3152), .IN3(n6290), .IN4(n5484), .Q(n3151)
         );
  OA22X1 U3701 ( .IN1(n6290), .IN2(n5475), .IN3(n5273), .IN4(n6136), .Q(n3152)
         );
  OAI22X1 U3702 ( .IN1(n6445), .IN2(n5526), .IN3(n5521), .IN4(n3153), .QN(
        N10494) );
  OA22X1 U3703 ( .IN1(n6445), .IN2(n5498), .IN3(n5505), .IN4(n3154), .Q(n3153)
         );
  OA22X1 U3704 ( .IN1(n5488), .IN2(n3155), .IN3(n6291), .IN4(n5484), .Q(n3154)
         );
  OA22X1 U3705 ( .IN1(n6291), .IN2(n5474), .IN3(n5273), .IN4(n6137), .Q(n3155)
         );
  OAI22X1 U3706 ( .IN1(n6446), .IN2(n5527), .IN3(n5521), .IN4(n3156), .QN(
        N10493) );
  OA22X1 U3707 ( .IN1(n6446), .IN2(n5498), .IN3(n5506), .IN4(n3157), .Q(n3156)
         );
  OA22X1 U3708 ( .IN1(n5488), .IN2(n3158), .IN3(n6292), .IN4(n5484), .Q(n3157)
         );
  OA22X1 U3709 ( .IN1(n6292), .IN2(n5476), .IN3(n5273), .IN4(n6138), .Q(n3158)
         );
  OAI22X1 U3710 ( .IN1(n6447), .IN2(n5516), .IN3(n5521), .IN4(n3159), .QN(
        N10492) );
  OA22X1 U3711 ( .IN1(n6447), .IN2(n5498), .IN3(n5506), .IN4(n3160), .Q(n3159)
         );
  OA22X1 U3712 ( .IN1(n5488), .IN2(n3161), .IN3(n6293), .IN4(n5484), .Q(n3160)
         );
  OA22X1 U3713 ( .IN1(n6293), .IN2(n5478), .IN3(n5273), .IN4(n6139), .Q(n3161)
         );
  OAI22X1 U3714 ( .IN1(n6448), .IN2(n5516), .IN3(n5521), .IN4(n3162), .QN(
        N10491) );
  OA22X1 U3715 ( .IN1(n6448), .IN2(n5498), .IN3(n5506), .IN4(n3163), .Q(n3162)
         );
  OA22X1 U3716 ( .IN1(n5487), .IN2(n3164), .IN3(n6294), .IN4(n5484), .Q(n3163)
         );
  OA22X1 U3717 ( .IN1(n6294), .IN2(n5480), .IN3(n5273), .IN4(n6140), .Q(n3164)
         );
  OAI22X1 U3718 ( .IN1(n6449), .IN2(n5522), .IN3(n5521), .IN4(n3165), .QN(
        N10490) );
  OA22X1 U3719 ( .IN1(n6449), .IN2(n5498), .IN3(n5506), .IN4(n3166), .Q(n3165)
         );
  OA22X1 U3720 ( .IN1(n5487), .IN2(n3167), .IN3(n6295), .IN4(n5484), .Q(n3166)
         );
  OA22X1 U3721 ( .IN1(n6295), .IN2(n5478), .IN3(n5273), .IN4(n6141), .Q(n3167)
         );
  OAI22X1 U3722 ( .IN1(n6450), .IN2(n5523), .IN3(n5521), .IN4(n3168), .QN(
        N10489) );
  OA22X1 U3723 ( .IN1(n6450), .IN2(n5498), .IN3(n5506), .IN4(n3169), .Q(n3168)
         );
  OA22X1 U3724 ( .IN1(n5487), .IN2(n3170), .IN3(n6296), .IN4(n5484), .Q(n3169)
         );
  OA22X1 U3725 ( .IN1(n6296), .IN2(n5473), .IN3(n5273), .IN4(n6142), .Q(n3170)
         );
  OAI22X1 U3726 ( .IN1(n6451), .IN2(n5524), .IN3(n5521), .IN4(n3171), .QN(
        N10488) );
  OA22X1 U3727 ( .IN1(n6451), .IN2(n5497), .IN3(n5507), .IN4(n3172), .Q(n3171)
         );
  OA22X1 U3728 ( .IN1(n5487), .IN2(n3173), .IN3(n6297), .IN4(n5484), .Q(n3172)
         );
  OA22X1 U3729 ( .IN1(n6297), .IN2(n5474), .IN3(n5273), .IN4(n6143), .Q(n3173)
         );
  OAI22X1 U3730 ( .IN1(n6452), .IN2(n5525), .IN3(n5521), .IN4(n3174), .QN(
        N10487) );
  OA22X1 U3731 ( .IN1(n6452), .IN2(n5497), .IN3(n5507), .IN4(n3175), .Q(n3174)
         );
  OA22X1 U3732 ( .IN1(n5487), .IN2(n3176), .IN3(n6298), .IN4(n5484), .Q(n3175)
         );
  OA22X1 U3733 ( .IN1(n6298), .IN2(n5479), .IN3(n5273), .IN4(n6144), .Q(n3176)
         );
  OAI22X1 U3734 ( .IN1(n6453), .IN2(n5526), .IN3(n5521), .IN4(n3177), .QN(
        N10486) );
  OA22X1 U3735 ( .IN1(n6453), .IN2(n5497), .IN3(n5507), .IN4(n3178), .Q(n3177)
         );
  OA22X1 U3736 ( .IN1(n5487), .IN2(n3179), .IN3(n6299), .IN4(n5484), .Q(n3178)
         );
  OA22X1 U3737 ( .IN1(n6299), .IN2(n5477), .IN3(n5273), .IN4(n6145), .Q(n3179)
         );
  OAI22X1 U3738 ( .IN1(n6454), .IN2(n5527), .IN3(n5518), .IN4(n3180), .QN(
        N10485) );
  OA22X1 U3739 ( .IN1(n6454), .IN2(n5497), .IN3(n5507), .IN4(n3181), .Q(n3180)
         );
  OA22X1 U3740 ( .IN1(n5487), .IN2(n3182), .IN3(n6300), .IN4(n5484), .Q(n3181)
         );
  OA22X1 U3741 ( .IN1(n6300), .IN2(n5475), .IN3(n5273), .IN4(n6146), .Q(n3182)
         );
  OA22X1 U3743 ( .IN1(n6320), .IN2(n5497), .IN3(n5507), .IN4(n3184), .Q(n3183)
         );
  OA22X1 U3747 ( .IN1(n6321), .IN2(n5497), .IN3(n5508), .IN4(n3187), .Q(n3186)
         );
  OA22X1 U3751 ( .IN1(n6322), .IN2(n5497), .IN3(n5508), .IN4(n3190), .Q(n3189)
         );
  OA22X1 U3755 ( .IN1(n6323), .IN2(n5497), .IN3(n5508), .IN4(n3193), .Q(n3192)
         );
  OA22X1 U3759 ( .IN1(n6324), .IN2(n5497), .IN3(n5508), .IN4(n3196), .Q(n3195)
         );
  OA22X1 U3763 ( .IN1(n6325), .IN2(n5497), .IN3(n5508), .IN4(n3199), .Q(n3198)
         );
  OA22X1 U3767 ( .IN1(n6326), .IN2(n5497), .IN3(n5509), .IN4(n3202), .Q(n3201)
         );
  OA22X1 U3771 ( .IN1(n6327), .IN2(n5497), .IN3(n5509), .IN4(n3205), .Q(n3204)
         );
  OA22X1 U3775 ( .IN1(n6328), .IN2(n5497), .IN3(n5509), .IN4(n3208), .Q(n3207)
         );
  OA22X1 U3779 ( .IN1(n6329), .IN2(n5497), .IN3(n5509), .IN4(n3211), .Q(n3210)
         );
  OA22X1 U3783 ( .IN1(n6330), .IN2(n5496), .IN3(n5509), .IN4(n3214), .Q(n3213)
         );
  OA22X1 U3787 ( .IN1(n6331), .IN2(n5496), .IN3(n5510), .IN4(n3217), .Q(n3216)
         );
  OA22X1 U3791 ( .IN1(n6332), .IN2(n5496), .IN3(n5510), .IN4(n3220), .Q(n3219)
         );
  OA22X1 U3795 ( .IN1(n6333), .IN2(n5496), .IN3(n5510), .IN4(n3223), .Q(n3222)
         );
  OA22X1 U3799 ( .IN1(n6334), .IN2(n5496), .IN3(n5510), .IN4(n3226), .Q(n3225)
         );
  OA22X1 U3803 ( .IN1(n6335), .IN2(n5496), .IN3(n5510), .IN4(n3229), .Q(n3228)
         );
  OA22X1 U3807 ( .IN1(n6336), .IN2(n5496), .IN3(n5511), .IN4(n3232), .Q(n3231)
         );
  OA22X1 U3811 ( .IN1(n6337), .IN2(n5496), .IN3(n5511), .IN4(n3235), .Q(n3234)
         );
  OA22X1 U3815 ( .IN1(n6338), .IN2(n5496), .IN3(n5511), .IN4(n3238), .Q(n3237)
         );
  OA22X1 U3819 ( .IN1(n6339), .IN2(n5496), .IN3(n5511), .IN4(n3241), .Q(n3240)
         );
  OA22X1 U3823 ( .IN1(n6340), .IN2(n5496), .IN3(n5511), .IN4(n3244), .Q(n3243)
         );
  OA22X1 U3827 ( .IN1(n6341), .IN2(n5496), .IN3(n5507), .IN4(n3247), .Q(n3246)
         );
  OA22X1 U3831 ( .IN1(n6342), .IN2(n5496), .IN3(n5512), .IN4(n3250), .Q(n3249)
         );
  OA22X1 U3835 ( .IN1(n6343), .IN2(n5496), .IN3(n5513), .IN4(n3253), .Q(n3252)
         );
  OA22X1 U3839 ( .IN1(n6344), .IN2(n5495), .IN3(n5509), .IN4(n3256), .Q(n3255)
         );
  OA22X1 U3843 ( .IN1(n6345), .IN2(n5495), .IN3(n5506), .IN4(n3259), .Q(n3258)
         );
  OA22X1 U3847 ( .IN1(n6346), .IN2(n5495), .IN3(n5508), .IN4(n3262), .Q(n3261)
         );
  OA22X1 U3851 ( .IN1(n6315), .IN2(n5495), .IN3(n5509), .IN4(n3265), .Q(n3264)
         );
  OA22X1 U3855 ( .IN1(n6316), .IN2(n5495), .IN3(n5504), .IN4(n3268), .Q(n3267)
         );
  OA22X1 U3859 ( .IN1(n6317), .IN2(n5495), .IN3(n5505), .IN4(n3271), .Q(n3270)
         );
  OA22X1 U3863 ( .IN1(n6318), .IN2(n5495), .IN3(n5506), .IN4(n3274), .Q(n3273)
         );
  OA22X1 U3867 ( .IN1(n6319), .IN2(n5495), .IN3(n5511), .IN4(n3277), .Q(n3276)
         );
  OAI22X1 U3870 ( .IN1(n6455), .IN2(n5522), .IN3(n5517), .IN4(n3279), .QN(
        N10452) );
  OA22X1 U3871 ( .IN1(n6455), .IN2(n5495), .IN3(n5510), .IN4(n3280), .Q(n3279)
         );
  OA22X1 U3872 ( .IN1(n5487), .IN2(n3281), .IN3(n6301), .IN4(n5483), .Q(n3280)
         );
  OA22X1 U3873 ( .IN1(n6301), .IN2(n5476), .IN3(n5273), .IN4(n6147), .Q(n3281)
         );
  OAI22X1 U3874 ( .IN1(n6456), .IN2(n5525), .IN3(n5518), .IN4(n3282), .QN(
        N10451) );
  OA22X1 U3875 ( .IN1(n6456), .IN2(n5495), .IN3(n5508), .IN4(n3283), .Q(n3282)
         );
  OA22X1 U3876 ( .IN1(n5487), .IN2(n3284), .IN3(n6302), .IN4(n5483), .Q(n3283)
         );
  OA22X1 U3877 ( .IN1(n6302), .IN2(n5477), .IN3(n5273), .IN4(n6148), .Q(n3284)
         );
  OAI22X1 U3878 ( .IN1(n6457), .IN2(n5526), .IN3(n5517), .IN4(n3285), .QN(
        N10450) );
  OA22X1 U3879 ( .IN1(n6457), .IN2(n5495), .IN3(n5508), .IN4(n3286), .Q(n3285)
         );
  OA22X1 U3880 ( .IN1(n5487), .IN2(n3287), .IN3(n6303), .IN4(n5483), .Q(n3286)
         );
  OA22X1 U3881 ( .IN1(n6303), .IN2(n5479), .IN3(n5273), .IN4(n6149), .Q(n3287)
         );
  OAI22X1 U3882 ( .IN1(n6458), .IN2(n5527), .IN3(n5518), .IN4(n3288), .QN(
        N10449) );
  OA22X1 U3883 ( .IN1(n6458), .IN2(n5495), .IN3(n5512), .IN4(n3289), .Q(n3288)
         );
  OA22X1 U3884 ( .IN1(n5487), .IN2(n3290), .IN3(n6304), .IN4(n5483), .Q(n3289)
         );
  OA22X1 U3885 ( .IN1(n6304), .IN2(n5474), .IN3(n5273), .IN4(n6150), .Q(n3290)
         );
  OAI22X1 U3886 ( .IN1(n6459), .IN2(n5516), .IN3(n5517), .IN4(n3291), .QN(
        N10448) );
  OA22X1 U3887 ( .IN1(n6459), .IN2(n5495), .IN3(n5512), .IN4(n3292), .Q(n3291)
         );
  OA22X1 U3888 ( .IN1(n5487), .IN2(n3293), .IN3(n6305), .IN4(n5483), .Q(n3292)
         );
  OA22X1 U3889 ( .IN1(n6305), .IN2(n5480), .IN3(n5471), .IN4(n6151), .Q(n3293)
         );
  NAND4X0 U3890 ( .IN1(n3294), .IN2(n5495), .IN3(n3295), .IN4(n5483), .QN(
        decodedVector_o[6]) );
  NAND4X0 U3892 ( .IN1(decodedPacketValid[4]), .IN2(N2173), .IN3(n2908), .IN4(
        n5995), .QN(n2918) );
  NAND4X0 U3893 ( .IN1(decodedPacketValid[7]), .IN2(N8581), .IN3(n2909), .IN4(
        n5992), .QN(n2912) );
  NAND4X0 U3894 ( .IN1(decodedPacketValid[6]), .IN2(N6445), .IN3(n2910), .IN4(
        n5993), .QN(n2914) );
  NAND4X0 U3895 ( .IN1(decodedPacketValid[3]), .IN2(N1069), .IN3(N1070), .IN4(
        n5996), .QN(n3294) );
  OA22X1 U3913 ( .IN1(n5856), .IN2(n5444), .IN3(n5448), .IN4(n3313), .Q(n3312)
         );
  OAI22X1 U3916 ( .IN1(n6384), .IN2(n5468), .IN3(n5460), .IN4(n3315), .QN(
        N10441) );
  OA22X1 U3917 ( .IN1(n6349), .IN2(n5444), .IN3(n5454), .IN4(n3316), .Q(n3315)
         );
  OA22X1 U3918 ( .IN1(n5435), .IN2(n3317), .IN3(n6230), .IN4(n5427), .Q(n3316)
         );
  OA22X1 U3919 ( .IN1(n6195), .IN2(n5414), .IN3(n5271), .IN4(n6076), .Q(n3317)
         );
  OAI22X1 U3920 ( .IN1(n6376), .IN2(n5468), .IN3(n5460), .IN4(n3318), .QN(
        N10440) );
  OA22X1 U3921 ( .IN1(n6348), .IN2(n5444), .IN3(n5448), .IN4(n3319), .Q(n3318)
         );
  OA22X1 U3922 ( .IN1(n5435), .IN2(n3320), .IN3(n6222), .IN4(n5427), .Q(n3319)
         );
  OA22X1 U3923 ( .IN1(n6194), .IN2(n5414), .IN3(n5413), .IN4(n6068), .Q(n3320)
         );
  OAI22X1 U3924 ( .IN1(n6373), .IN2(n5468), .IN3(n5460), .IN4(n3321), .QN(
        N10439) );
  OA22X1 U3925 ( .IN1(n6374), .IN2(n5444), .IN3(n5445), .IN4(n3322), .Q(n3321)
         );
  OA22X1 U3926 ( .IN1(n5435), .IN2(n3323), .IN3(n6219), .IN4(n5427), .Q(n3322)
         );
  OA22X1 U3927 ( .IN1(n6220), .IN2(n5414), .IN3(n5413), .IN4(n6064), .Q(n3323)
         );
  OA22X1 U3929 ( .IN1(n6371), .IN2(n5444), .IN3(n5452), .IN4(n3325), .Q(n3324)
         );
  OAI22X1 U3932 ( .IN1(n6373), .IN2(n5468), .IN3(n5460), .IN4(n3327), .QN(
        N10437) );
  OA22X1 U3933 ( .IN1(n6370), .IN2(n5444), .IN3(n5451), .IN4(n3328), .Q(n3327)
         );
  OA22X1 U3934 ( .IN1(n5435), .IN2(n3329), .IN3(n6219), .IN4(n5427), .Q(n3328)
         );
  OA22X1 U3935 ( .IN1(n6216), .IN2(n5414), .IN3(n5413), .IN4(n6065), .Q(n3329)
         );
  OAI22X1 U3936 ( .IN1(n6395), .IN2(n5468), .IN3(n5461), .IN4(n3330), .QN(
        N10436) );
  OA22X1 U3937 ( .IN1(n6347), .IN2(n5444), .IN3(n5450), .IN4(n3331), .Q(n3330)
         );
  OA22X1 U3938 ( .IN1(n5434), .IN2(n3332), .IN3(n6245), .IN4(n5427), .Q(n3331)
         );
  OA22X1 U3939 ( .IN1(n6193), .IN2(n5414), .IN3(n5413), .IN4(n6091), .Q(n3332)
         );
  OAI22X1 U3940 ( .IN1(n5967), .IN2(n5468), .IN3(n5461), .IN4(n3333), .QN(
        N10435) );
  OA22X1 U3941 ( .IN1(n6369), .IN2(n5444), .IN3(n5445), .IN4(n3334), .Q(n3333)
         );
  OA22X1 U3942 ( .IN1(n5434), .IN2(n3335), .IN3(n5952), .IN4(n5427), .Q(n3334)
         );
  OA22X1 U3943 ( .IN1(n6215), .IN2(n5415), .IN3(n5413), .IN4(n5937), .Q(n3335)
         );
  OAI22X1 U3944 ( .IN1(n5968), .IN2(n5467), .IN3(n5461), .IN4(n3336), .QN(
        N10434) );
  OA22X1 U3945 ( .IN1(n6368), .IN2(n5444), .IN3(n5446), .IN4(n3337), .Q(n3336)
         );
  OA22X1 U3946 ( .IN1(n5434), .IN2(n3338), .IN3(n5953), .IN4(n5427), .Q(n3337)
         );
  OA22X1 U3947 ( .IN1(n6214), .IN2(n5415), .IN3(n5413), .IN4(n5938), .Q(n3338)
         );
  OAI22X1 U3948 ( .IN1(n5969), .IN2(n5467), .IN3(n5461), .IN4(n3339), .QN(
        N10433) );
  OA22X1 U3949 ( .IN1(n6367), .IN2(n5444), .IN3(n5447), .IN4(n3340), .Q(n3339)
         );
  OA22X1 U3950 ( .IN1(n5434), .IN2(n3341), .IN3(n5954), .IN4(n5427), .Q(n3340)
         );
  OA22X1 U3951 ( .IN1(n6213), .IN2(n5415), .IN3(n5413), .IN4(n5939), .Q(n3341)
         );
  OAI22X1 U3952 ( .IN1(n5970), .IN2(n5467), .IN3(n5461), .IN4(n3342), .QN(
        N10432) );
  OA22X1 U3953 ( .IN1(n6366), .IN2(n5444), .IN3(n5455), .IN4(n3343), .Q(n3342)
         );
  OA22X1 U3954 ( .IN1(n5434), .IN2(n3344), .IN3(n5955), .IN4(n5427), .Q(n3343)
         );
  OA22X1 U3955 ( .IN1(n6212), .IN2(n5415), .IN3(n5413), .IN4(n5940), .Q(n3344)
         );
  OAI22X1 U3956 ( .IN1(n5971), .IN2(n5467), .IN3(n5461), .IN4(n3345), .QN(
        N10431) );
  OA22X1 U3957 ( .IN1(n6365), .IN2(n5443), .IN3(n5449), .IN4(n3346), .Q(n3345)
         );
  OA22X1 U3958 ( .IN1(n5434), .IN2(n3347), .IN3(n5956), .IN4(n5427), .Q(n3346)
         );
  OA22X1 U3959 ( .IN1(n6211), .IN2(n5415), .IN3(n5413), .IN4(n5941), .Q(n3347)
         );
  OAI22X1 U3960 ( .IN1(n5972), .IN2(n5467), .IN3(n5461), .IN4(n3348), .QN(
        N10430) );
  OA22X1 U3961 ( .IN1(n6364), .IN2(n5443), .IN3(n5452), .IN4(n3349), .Q(n3348)
         );
  OA22X1 U3962 ( .IN1(n5434), .IN2(n3350), .IN3(n5957), .IN4(n5427), .Q(n3349)
         );
  OA22X1 U3963 ( .IN1(n6210), .IN2(n5418), .IN3(n5413), .IN4(n5942), .Q(n3350)
         );
  OAI22X1 U3964 ( .IN1(n5973), .IN2(n5467), .IN3(n5461), .IN4(n3351), .QN(
        N10429) );
  OA22X1 U3965 ( .IN1(n6363), .IN2(n5443), .IN3(n5451), .IN4(n3352), .Q(n3351)
         );
  OA22X1 U3966 ( .IN1(n5434), .IN2(n3353), .IN3(n5958), .IN4(n5427), .Q(n3352)
         );
  OA22X1 U3967 ( .IN1(n6209), .IN2(n5415), .IN3(n5413), .IN4(n5943), .Q(n3353)
         );
  OAI22X1 U3968 ( .IN1(n5974), .IN2(n5467), .IN3(n5461), .IN4(n3354), .QN(
        N10428) );
  OA22X1 U3969 ( .IN1(n6362), .IN2(n5443), .IN3(n5455), .IN4(n3355), .Q(n3354)
         );
  OA22X1 U3970 ( .IN1(n5434), .IN2(n3356), .IN3(n5959), .IN4(n5427), .Q(n3355)
         );
  OA22X1 U3971 ( .IN1(n6208), .IN2(n5417), .IN3(n5413), .IN4(n5944), .Q(n3356)
         );
  OAI22X1 U3972 ( .IN1(n5975), .IN2(n5466), .IN3(n5461), .IN4(n3357), .QN(
        N10427) );
  OA22X1 U3973 ( .IN1(n6308), .IN2(n5443), .IN3(n5454), .IN4(n3358), .Q(n3357)
         );
  OA22X1 U3974 ( .IN1(n5434), .IN2(n3359), .IN3(n5960), .IN4(n5426), .Q(n3358)
         );
  OA22X1 U3975 ( .IN1(n6154), .IN2(n5419), .IN3(n5413), .IN4(n5945), .Q(n3359)
         );
  OAI22X1 U3976 ( .IN1(n5976), .IN2(n5466), .IN3(n5461), .IN4(n3360), .QN(
        N10426) );
  OA22X1 U3977 ( .IN1(n6309), .IN2(n5443), .IN3(n5445), .IN4(n3361), .Q(n3360)
         );
  OA22X1 U3978 ( .IN1(n5434), .IN2(n3362), .IN3(n5961), .IN4(n5426), .Q(n3361)
         );
  OA22X1 U3979 ( .IN1(n6155), .IN2(n5420), .IN3(n5413), .IN4(n5946), .Q(n3362)
         );
  OAI22X1 U3980 ( .IN1(n5977), .IN2(n5466), .IN3(n5461), .IN4(n3363), .QN(
        N10425) );
  OA22X1 U3981 ( .IN1(n6310), .IN2(n5443), .IN3(n5448), .IN4(n3364), .Q(n3363)
         );
  OA22X1 U3982 ( .IN1(n5434), .IN2(n3365), .IN3(n5962), .IN4(n5426), .Q(n3364)
         );
  OA22X1 U3983 ( .IN1(n6156), .IN2(n5417), .IN3(n5413), .IN4(n5947), .Q(n3365)
         );
  OAI22X1 U3984 ( .IN1(n5978), .IN2(n5466), .IN3(n5461), .IN4(n3366), .QN(
        N10424) );
  OA22X1 U3985 ( .IN1(n6311), .IN2(n5443), .IN3(n5455), .IN4(n3367), .Q(n3366)
         );
  OA22X1 U3986 ( .IN1(n5433), .IN2(n3368), .IN3(n5963), .IN4(n5426), .Q(n3367)
         );
  OA22X1 U3987 ( .IN1(n6157), .IN2(n5415), .IN3(n5413), .IN4(n5948), .Q(n3368)
         );
  OAI22X1 U3988 ( .IN1(n5979), .IN2(n5466), .IN3(n5461), .IN4(n3369), .QN(
        N10423) );
  OA22X1 U3989 ( .IN1(n6312), .IN2(n5443), .IN3(n5454), .IN4(n3370), .Q(n3369)
         );
  OA22X1 U3990 ( .IN1(n5433), .IN2(n3371), .IN3(n5964), .IN4(n5426), .Q(n3370)
         );
  OA22X1 U3991 ( .IN1(n6158), .IN2(n5417), .IN3(n5413), .IN4(n5949), .Q(n3371)
         );
  OAI22X1 U3992 ( .IN1(n5980), .IN2(n5466), .IN3(n5461), .IN4(n3372), .QN(
        N10422) );
  OA22X1 U3993 ( .IN1(n6313), .IN2(n5443), .IN3(n5453), .IN4(n3373), .Q(n3372)
         );
  OA22X1 U3994 ( .IN1(n5433), .IN2(n3374), .IN3(n5965), .IN4(n5426), .Q(n3373)
         );
  OA22X1 U3995 ( .IN1(n6159), .IN2(n5416), .IN3(n5413), .IN4(n5950), .Q(n3374)
         );
  OAI22X1 U3996 ( .IN1(n5981), .IN2(n5466), .IN3(n5461), .IN4(n3375), .QN(
        N10421) );
  OA22X1 U3997 ( .IN1(n6314), .IN2(n5443), .IN3(n5454), .IN4(n3376), .Q(n3375)
         );
  OA22X1 U3998 ( .IN1(n5433), .IN2(n3377), .IN3(n5966), .IN4(n5426), .Q(n3376)
         );
  OA22X1 U3999 ( .IN1(n6160), .IN2(n5414), .IN3(n5413), .IN4(n5951), .Q(n3377)
         );
  OAI22X1 U4000 ( .IN1(n6375), .IN2(n5468), .IN3(n5461), .IN4(n3378), .QN(
        N10420) );
  OA22X1 U4001 ( .IN1(n6307), .IN2(n5443), .IN3(n5453), .IN4(n3379), .Q(n3378)
         );
  OA22X1 U4002 ( .IN1(n5433), .IN2(n3380), .IN3(n6221), .IN4(n5426), .Q(n3379)
         );
  OA22X1 U4003 ( .IN1(n6153), .IN2(n5416), .IN3(n5413), .IN4(n6067), .Q(n3380)
         );
  OAI22X1 U4004 ( .IN1(n6372), .IN2(n5457), .IN3(n5461), .IN4(n3381), .QN(
        N10418) );
  OA22X1 U4005 ( .IN1(n6306), .IN2(n5443), .IN3(n5454), .IN4(n3382), .Q(n3381)
         );
  OA22X1 U4006 ( .IN1(n5433), .IN2(n3383), .IN3(n6218), .IN4(n5426), .Q(n3382)
         );
  OA22X1 U4007 ( .IN1(n6152), .IN2(n5416), .IN3(n5413), .IN4(n6064), .Q(n3383)
         );
  OAI22X1 U4008 ( .IN1(n6377), .IN2(n5456), .IN3(n5461), .IN4(n3384), .QN(
        N10416) );
  OA22X1 U4009 ( .IN1(n6422), .IN2(n5443), .IN3(n5455), .IN4(n3385), .Q(n3384)
         );
  OA22X1 U4010 ( .IN1(n5433), .IN2(n3386), .IN3(n6223), .IN4(n5426), .Q(n3385)
         );
  OA22X1 U4011 ( .IN1(n6268), .IN2(n5416), .IN3(n5413), .IN4(n6069), .Q(n3386)
         );
  OAI22X1 U4012 ( .IN1(n6378), .IN2(n5463), .IN3(n5461), .IN4(n3387), .QN(
        N10415) );
  OA22X1 U4013 ( .IN1(n6421), .IN2(n5442), .IN3(n5451), .IN4(n3388), .Q(n3387)
         );
  OA22X1 U4014 ( .IN1(n5433), .IN2(n3389), .IN3(n6224), .IN4(n5426), .Q(n3388)
         );
  OA22X1 U4015 ( .IN1(n6267), .IN2(n5416), .IN3(n5413), .IN4(n6070), .Q(n3389)
         );
  OAI22X1 U4016 ( .IN1(n6379), .IN2(n5465), .IN3(n5461), .IN4(n3390), .QN(
        N10414) );
  OA22X1 U4017 ( .IN1(n6420), .IN2(n5442), .IN3(n5448), .IN4(n3391), .Q(n3390)
         );
  OA22X1 U4018 ( .IN1(n5433), .IN2(n3392), .IN3(n6225), .IN4(n5426), .Q(n3391)
         );
  OA22X1 U4019 ( .IN1(n6266), .IN2(n5416), .IN3(n5413), .IN4(n6071), .Q(n3392)
         );
  OAI22X1 U4020 ( .IN1(n6380), .IN2(n5463), .IN3(n5461), .IN4(n3393), .QN(
        N10413) );
  OA22X1 U4021 ( .IN1(n6419), .IN2(n5442), .IN3(n5453), .IN4(n3394), .Q(n3393)
         );
  OA22X1 U4022 ( .IN1(n5433), .IN2(n3395), .IN3(n6226), .IN4(n5426), .Q(n3394)
         );
  OA22X1 U4023 ( .IN1(n6265), .IN2(n5417), .IN3(n5413), .IN4(n6072), .Q(n3395)
         );
  OAI22X1 U4024 ( .IN1(n6381), .IN2(n5464), .IN3(n5461), .IN4(n3396), .QN(
        N10412) );
  OA22X1 U4025 ( .IN1(n6418), .IN2(n5442), .IN3(n5453), .IN4(n3397), .Q(n3396)
         );
  OA22X1 U4026 ( .IN1(n5433), .IN2(n3398), .IN3(n6227), .IN4(n5426), .Q(n3397)
         );
  OA22X1 U4027 ( .IN1(n6264), .IN2(n5417), .IN3(n5413), .IN4(n6073), .Q(n3398)
         );
  OAI22X1 U4028 ( .IN1(n6382), .IN2(n5468), .IN3(n5461), .IN4(n3399), .QN(
        N10411) );
  OA22X1 U4029 ( .IN1(n6417), .IN2(n5442), .IN3(n5454), .IN4(n3400), .Q(n3399)
         );
  OA22X1 U4030 ( .IN1(n5433), .IN2(n3401), .IN3(n6228), .IN4(n5426), .Q(n3400)
         );
  OA22X1 U4031 ( .IN1(n6263), .IN2(n5417), .IN3(n5413), .IN4(n6074), .Q(n3401)
         );
  OAI22X1 U4032 ( .IN1(n6383), .IN2(n5466), .IN3(n5461), .IN4(n3402), .QN(
        N10410) );
  OA22X1 U4033 ( .IN1(n6416), .IN2(n5442), .IN3(n5455), .IN4(n3403), .Q(n3402)
         );
  OA22X1 U4034 ( .IN1(n5432), .IN2(n3404), .IN3(n6229), .IN4(n5426), .Q(n3403)
         );
  OA22X1 U4035 ( .IN1(n6262), .IN2(n5417), .IN3(n5413), .IN4(n6075), .Q(n3404)
         );
  OAI22X1 U4036 ( .IN1(n6385), .IN2(n5467), .IN3(n5461), .IN4(n3405), .QN(
        N10409) );
  OA22X1 U4037 ( .IN1(n6359), .IN2(n5442), .IN3(n5452), .IN4(n3406), .Q(n3405)
         );
  OA22X1 U4038 ( .IN1(n5432), .IN2(n3407), .IN3(n6231), .IN4(n5426), .Q(n3406)
         );
  OA22X1 U4039 ( .IN1(n6205), .IN2(n5417), .IN3(n5413), .IN4(n6077), .Q(n3407)
         );
  OAI22X1 U4040 ( .IN1(n6386), .IN2(n5457), .IN3(n5461), .IN4(n3408), .QN(
        N10408) );
  OA22X1 U4041 ( .IN1(n6358), .IN2(n5442), .IN3(n5446), .IN4(n3409), .Q(n3408)
         );
  OA22X1 U4042 ( .IN1(n5432), .IN2(n3410), .IN3(n6232), .IN4(n5426), .Q(n3409)
         );
  OA22X1 U4043 ( .IN1(n6204), .IN2(n5418), .IN3(n5413), .IN4(n6078), .Q(n3410)
         );
  OAI22X1 U4044 ( .IN1(n6387), .IN2(n5456), .IN3(n5461), .IN4(n3411), .QN(
        N10407) );
  OA22X1 U4045 ( .IN1(n6357), .IN2(n5442), .IN3(n5448), .IN4(n3412), .Q(n3411)
         );
  OA22X1 U4046 ( .IN1(n5432), .IN2(n3413), .IN3(n6233), .IN4(n5426), .Q(n3412)
         );
  OA22X1 U4047 ( .IN1(n6203), .IN2(n5414), .IN3(n5413), .IN4(n6079), .Q(n3413)
         );
  OAI22X1 U4048 ( .IN1(n6388), .IN2(n5463), .IN3(n5461), .IN4(n3414), .QN(
        N10406) );
  OA22X1 U4049 ( .IN1(n6356), .IN2(n5442), .IN3(n5452), .IN4(n3415), .Q(n3414)
         );
  OA22X1 U4050 ( .IN1(n5432), .IN2(n3416), .IN3(n6234), .IN4(n5426), .Q(n3415)
         );
  OA22X1 U4051 ( .IN1(n6202), .IN2(n5416), .IN3(n5413), .IN4(n6080), .Q(n3416)
         );
  OAI22X1 U4052 ( .IN1(n6389), .IN2(n5465), .IN3(n5461), .IN4(n3417), .QN(
        N10405) );
  OA22X1 U4053 ( .IN1(n6355), .IN2(n5442), .IN3(n5451), .IN4(n3418), .Q(n3417)
         );
  OA22X1 U4054 ( .IN1(n5432), .IN2(n3419), .IN3(n6235), .IN4(n5426), .Q(n3418)
         );
  OA22X1 U4055 ( .IN1(n6201), .IN2(n5418), .IN3(n5412), .IN4(n6081), .Q(n3419)
         );
  OAI22X1 U4056 ( .IN1(n6390), .IN2(n5456), .IN3(n5461), .IN4(n3420), .QN(
        N10404) );
  OA22X1 U4057 ( .IN1(n6354), .IN2(n5442), .IN3(n5449), .IN4(n3421), .Q(n3420)
         );
  OA22X1 U4058 ( .IN1(n5432), .IN2(n3422), .IN3(n6236), .IN4(n5426), .Q(n3421)
         );
  OA22X1 U4059 ( .IN1(n6200), .IN2(n5419), .IN3(n5412), .IN4(n6082), .Q(n3422)
         );
  OAI22X1 U4060 ( .IN1(n6391), .IN2(n5463), .IN3(n5461), .IN4(n3423), .QN(
        N10403) );
  OA22X1 U4061 ( .IN1(n6353), .IN2(n5442), .IN3(n5450), .IN4(n3424), .Q(n3423)
         );
  OA22X1 U4062 ( .IN1(n5432), .IN2(n3425), .IN3(n6237), .IN4(n5426), .Q(n3424)
         );
  OA22X1 U4063 ( .IN1(n6199), .IN2(n5419), .IN3(n5412), .IN4(n6083), .Q(n3425)
         );
  OAI22X1 U4064 ( .IN1(n6400), .IN2(n5464), .IN3(n5461), .IN4(n3426), .QN(
        N10402) );
  OA22X1 U4065 ( .IN1(n6415), .IN2(n5442), .IN3(n5445), .IN4(n3427), .Q(n3426)
         );
  OA22X1 U4066 ( .IN1(n5432), .IN2(n3428), .IN3(n6246), .IN4(n5426), .Q(n3427)
         );
  OA22X1 U4067 ( .IN1(n6261), .IN2(n5420), .IN3(n5412), .IN4(n6092), .Q(n3428)
         );
  OAI22X1 U4068 ( .IN1(n6406), .IN2(n5465), .IN3(n5461), .IN4(n3429), .QN(
        N10401) );
  OA22X1 U4069 ( .IN1(n6414), .IN2(n5441), .IN3(n5446), .IN4(n3430), .Q(n3429)
         );
  OA22X1 U4070 ( .IN1(n5432), .IN2(n3431), .IN3(n6252), .IN4(n5426), .Q(n3430)
         );
  OA22X1 U4071 ( .IN1(n6260), .IN2(n5421), .IN3(n5412), .IN4(n6098), .Q(n3431)
         );
  OAI22X1 U4072 ( .IN1(n6407), .IN2(n5468), .IN3(n5461), .IN4(n3432), .QN(
        N10400) );
  OA22X1 U4073 ( .IN1(n6413), .IN2(n5441), .IN3(n5447), .IN4(n3433), .Q(n3432)
         );
  OA22X1 U4074 ( .IN1(n5432), .IN2(n3434), .IN3(n6253), .IN4(n5426), .Q(n3433)
         );
  OA22X1 U4075 ( .IN1(n6259), .IN2(n5415), .IN3(n5412), .IN4(n6099), .Q(n3434)
         );
  OAI22X1 U4076 ( .IN1(n6408), .IN2(n5457), .IN3(n5461), .IN4(n3435), .QN(
        N10399) );
  OA22X1 U4077 ( .IN1(n6412), .IN2(n5441), .IN3(n5452), .IN4(n3436), .Q(n3435)
         );
  OA22X1 U4078 ( .IN1(n5432), .IN2(n3437), .IN3(n6254), .IN4(n5426), .Q(n3436)
         );
  OA22X1 U4079 ( .IN1(n6258), .IN2(n5414), .IN3(n5412), .IN4(n6100), .Q(n3437)
         );
  OAI22X1 U4080 ( .IN1(n6409), .IN2(n5456), .IN3(n5461), .IN4(n3438), .QN(
        N10398) );
  OA22X1 U4081 ( .IN1(n6411), .IN2(n5441), .IN3(n5446), .IN4(n3439), .Q(n3438)
         );
  OA22X1 U4082 ( .IN1(n5431), .IN2(n3440), .IN3(n6255), .IN4(n5426), .Q(n3439)
         );
  OA22X1 U4083 ( .IN1(n6257), .IN2(n5418), .IN3(n5412), .IN4(n6101), .Q(n3440)
         );
  OAI22X1 U4084 ( .IN1(n6401), .IN2(n5465), .IN3(n5461), .IN4(n3441), .QN(
        N10397) );
  OA22X1 U4085 ( .IN1(n6410), .IN2(n5441), .IN3(n5448), .IN4(n3442), .Q(n3441)
         );
  OA22X1 U4086 ( .IN1(n5431), .IN2(n3443), .IN3(n6247), .IN4(n5426), .Q(n3442)
         );
  OA22X1 U4087 ( .IN1(n6256), .IN2(n5418), .IN3(n5412), .IN4(n6093), .Q(n3443)
         );
  OAI22X1 U4088 ( .IN1(n6399), .IN2(n5465), .IN3(n5461), .IN4(n3444), .QN(
        N10396) );
  OA22X1 U4089 ( .IN1(n6352), .IN2(n5441), .IN3(n5451), .IN4(n3445), .Q(n3444)
         );
  OA22X1 U4090 ( .IN1(n5431), .IN2(n3446), .IN3(n6244), .IN4(n5426), .Q(n3445)
         );
  OA22X1 U4091 ( .IN1(n6198), .IN2(n5418), .IN3(n5412), .IN4(n6090), .Q(n3446)
         );
  OAI22X1 U4092 ( .IN1(n6398), .IN2(n5465), .IN3(n5462), .IN4(n3447), .QN(
        N10395) );
  OA22X1 U4093 ( .IN1(n6402), .IN2(n5441), .IN3(n5445), .IN4(n3448), .Q(n3447)
         );
  OA22X1 U4094 ( .IN1(n5431), .IN2(n3449), .IN3(n6243), .IN4(n5426), .Q(n3448)
         );
  OA22X1 U4095 ( .IN1(n6248), .IN2(n5418), .IN3(n5412), .IN4(n6089), .Q(n3449)
         );
  OAI22X1 U4096 ( .IN1(n6397), .IN2(n5465), .IN3(n5462), .IN4(n3450), .QN(
        N10394) );
  OA22X1 U4097 ( .IN1(n6403), .IN2(n5441), .IN3(n5447), .IN4(n3451), .Q(n3450)
         );
  OA22X1 U4098 ( .IN1(n5431), .IN2(n3452), .IN3(n6242), .IN4(n5426), .Q(n3451)
         );
  OA22X1 U4099 ( .IN1(n6249), .IN2(n5418), .IN3(n5412), .IN4(n6091), .Q(n3452)
         );
  OAI22X1 U4100 ( .IN1(n6396), .IN2(n5465), .IN3(n5462), .IN4(n3453), .QN(
        N10393) );
  OA22X1 U4101 ( .IN1(n6404), .IN2(n5441), .IN3(n5449), .IN4(n3454), .Q(n3453)
         );
  OA22X1 U4102 ( .IN1(n5431), .IN2(n3455), .IN3(n6241), .IN4(n5426), .Q(n3454)
         );
  OA22X1 U4103 ( .IN1(n6250), .IN2(n5419), .IN3(n5412), .IN4(n6088), .Q(n3455)
         );
  OAI22X1 U4104 ( .IN1(n6399), .IN2(n5465), .IN3(n5462), .IN4(n3456), .QN(
        N10392) );
  OA22X1 U4105 ( .IN1(n6405), .IN2(n5441), .IN3(n5446), .IN4(n3457), .Q(n3456)
         );
  OA22X1 U4106 ( .IN1(n5431), .IN2(n3458), .IN3(n6243), .IN4(n5426), .Q(n3457)
         );
  OA22X1 U4107 ( .IN1(n6251), .IN2(n5419), .IN3(n5412), .IN4(n6087), .Q(n3458)
         );
  OAI22X1 U4108 ( .IN1(n6394), .IN2(n5465), .IN3(n5462), .IN4(n3459), .QN(
        N10391) );
  OA22X1 U4109 ( .IN1(n6393), .IN2(n5441), .IN3(n5455), .IN4(n3460), .Q(n3459)
         );
  OA22X1 U4110 ( .IN1(n5431), .IN2(n3461), .IN3(n6240), .IN4(n5426), .Q(n3460)
         );
  OA22X1 U4111 ( .IN1(n6239), .IN2(n5419), .IN3(n5412), .IN4(n6086), .Q(n3461)
         );
  OAI22X1 U4112 ( .IN1(n6361), .IN2(n5464), .IN3(n5462), .IN4(n3462), .QN(
        N10390) );
  OA22X1 U4113 ( .IN1(n6360), .IN2(n5441), .IN3(n5451), .IN4(n3463), .Q(n3462)
         );
  OA22X1 U4114 ( .IN1(n5431), .IN2(n3464), .IN3(n6207), .IN4(n5425), .Q(n3463)
         );
  OA22X1 U4115 ( .IN1(n6206), .IN2(n5419), .IN3(n5412), .IN4(n6053), .Q(n3464)
         );
  OAI22X1 U4116 ( .IN1(n6350), .IN2(n5464), .IN3(n5462), .IN4(n3465), .QN(
        N10389) );
  OA22X1 U4117 ( .IN1(n6351), .IN2(n5441), .IN3(n5451), .IN4(n3466), .Q(n3465)
         );
  OA22X1 U4118 ( .IN1(n5431), .IN2(n3467), .IN3(n6196), .IN4(n5425), .Q(n3466)
         );
  OA22X1 U4119 ( .IN1(n6197), .IN2(n5419), .IN3(n5412), .IN4(n6042), .Q(n3467)
         );
  OAI22X1 U4120 ( .IN1(n6395), .IN2(n5464), .IN3(n5462), .IN4(n3468), .QN(
        N10388) );
  OA22X1 U4121 ( .IN1(n6392), .IN2(n5441), .IN3(n5452), .IN4(n3469), .Q(n3468)
         );
  OA22X1 U4122 ( .IN1(n5431), .IN2(n3470), .IN3(n6242), .IN4(n5425), .Q(n3469)
         );
  OA22X1 U4123 ( .IN1(n6238), .IN2(n5420), .IN3(n5412), .IN4(n6088), .Q(n3470)
         );
  OAI22X1 U4124 ( .IN1(n6423), .IN2(n5464), .IN3(n5462), .IN4(n3471), .QN(
        N10387) );
  OA22X1 U4125 ( .IN1(n6423), .IN2(n5440), .IN3(n5453), .IN4(n3472), .Q(n3471)
         );
  OA22X1 U4126 ( .IN1(n5431), .IN2(n3473), .IN3(n6269), .IN4(n5425), .Q(n3472)
         );
  OA22X1 U4127 ( .IN1(n6269), .IN2(n5420), .IN3(n5412), .IN4(n6115), .Q(n3473)
         );
  OAI22X1 U4128 ( .IN1(n6424), .IN2(n5464), .IN3(n5462), .IN4(n3474), .QN(
        N10386) );
  OA22X1 U4129 ( .IN1(n6424), .IN2(n5440), .IN3(n5448), .IN4(n3475), .Q(n3474)
         );
  OA22X1 U4130 ( .IN1(n5430), .IN2(n3476), .IN3(n6270), .IN4(n5425), .Q(n3475)
         );
  OA22X1 U4131 ( .IN1(n6270), .IN2(n5420), .IN3(n5412), .IN4(n6116), .Q(n3476)
         );
  OAI22X1 U4132 ( .IN1(n6425), .IN2(n5464), .IN3(n5462), .IN4(n3477), .QN(
        N10385) );
  OA22X1 U4133 ( .IN1(n6425), .IN2(n5440), .IN3(n5453), .IN4(n3478), .Q(n3477)
         );
  OA22X1 U4134 ( .IN1(n5430), .IN2(n3479), .IN3(n6271), .IN4(n5425), .Q(n3478)
         );
  OA22X1 U4135 ( .IN1(n6271), .IN2(n5420), .IN3(n5412), .IN4(n6117), .Q(n3479)
         );
  OAI22X1 U4136 ( .IN1(n6426), .IN2(n5464), .IN3(n5462), .IN4(n3480), .QN(
        N10384) );
  OA22X1 U4137 ( .IN1(n6426), .IN2(n5440), .IN3(n5448), .IN4(n3481), .Q(n3480)
         );
  OA22X1 U4138 ( .IN1(n5430), .IN2(n3482), .IN3(n6272), .IN4(n5425), .Q(n3481)
         );
  OA22X1 U4139 ( .IN1(n6272), .IN2(n5420), .IN3(n5412), .IN4(n6118), .Q(n3482)
         );
  OAI22X1 U4140 ( .IN1(n6427), .IN2(n5463), .IN3(n5462), .IN4(n3483), .QN(
        N10383) );
  OA22X1 U4141 ( .IN1(n6427), .IN2(n5440), .IN3(n5454), .IN4(n3484), .Q(n3483)
         );
  OA22X1 U4142 ( .IN1(n5430), .IN2(n3485), .IN3(n6273), .IN4(n5425), .Q(n3484)
         );
  OA22X1 U4143 ( .IN1(n6273), .IN2(n5421), .IN3(n5412), .IN4(n6119), .Q(n3485)
         );
  OAI22X1 U4144 ( .IN1(n6428), .IN2(n5457), .IN3(n5462), .IN4(n3486), .QN(
        N10382) );
  OA22X1 U4145 ( .IN1(n6428), .IN2(n5440), .IN3(n5453), .IN4(n3487), .Q(n3486)
         );
  OA22X1 U4146 ( .IN1(n5430), .IN2(n3488), .IN3(n6274), .IN4(n5425), .Q(n3487)
         );
  OA22X1 U4147 ( .IN1(n6274), .IN2(n5421), .IN3(n5412), .IN4(n6120), .Q(n3488)
         );
  OAI22X1 U4148 ( .IN1(n6429), .IN2(n5456), .IN3(n5462), .IN4(n3489), .QN(
        N10381) );
  OA22X1 U4149 ( .IN1(n6429), .IN2(n5440), .IN3(n5455), .IN4(n3490), .Q(n3489)
         );
  OA22X1 U4150 ( .IN1(n5430), .IN2(n3491), .IN3(n6275), .IN4(n5425), .Q(n3490)
         );
  OA22X1 U4151 ( .IN1(n6275), .IN2(n5421), .IN3(n5412), .IN4(n6121), .Q(n3491)
         );
  OAI22X1 U4152 ( .IN1(n6430), .IN2(n5468), .IN3(n5462), .IN4(n3492), .QN(
        N10380) );
  OA22X1 U4153 ( .IN1(n6430), .IN2(n5440), .IN3(n5450), .IN4(n3493), .Q(n3492)
         );
  OA22X1 U4154 ( .IN1(n5430), .IN2(n3494), .IN3(n6276), .IN4(n5425), .Q(n3493)
         );
  OA22X1 U4155 ( .IN1(n6276), .IN2(n5421), .IN3(n5412), .IN4(n6122), .Q(n3494)
         );
  OAI22X1 U4156 ( .IN1(n6431), .IN2(n5464), .IN3(n5462), .IN4(n3495), .QN(
        N10379) );
  OA22X1 U4157 ( .IN1(n6431), .IN2(n5440), .IN3(n5450), .IN4(n3496), .Q(n3495)
         );
  OA22X1 U4158 ( .IN1(n5430), .IN2(n3497), .IN3(n6277), .IN4(n5425), .Q(n3496)
         );
  OA22X1 U4159 ( .IN1(n6277), .IN2(n5421), .IN3(n5412), .IN4(n6123), .Q(n3497)
         );
  OAI22X1 U4160 ( .IN1(n6432), .IN2(n5466), .IN3(n5462), .IN4(n3498), .QN(
        N10378) );
  OA22X1 U4161 ( .IN1(n6432), .IN2(n5440), .IN3(n5447), .IN4(n3499), .Q(n3498)
         );
  OA22X1 U4162 ( .IN1(n5430), .IN2(n3500), .IN3(n6278), .IN4(n5425), .Q(n3499)
         );
  OA22X1 U4163 ( .IN1(n6278), .IN2(n5421), .IN3(n5412), .IN4(n6124), .Q(n3500)
         );
  OAI22X1 U4164 ( .IN1(n6433), .IN2(n5467), .IN3(n5462), .IN4(n3501), .QN(
        N10377) );
  OA22X1 U4165 ( .IN1(n6433), .IN2(n5440), .IN3(n5449), .IN4(n3502), .Q(n3501)
         );
  OA22X1 U4166 ( .IN1(n5430), .IN2(n3503), .IN3(n6279), .IN4(n5425), .Q(n3502)
         );
  OA22X1 U4167 ( .IN1(n6279), .IN2(n5416), .IN3(n5412), .IN4(n6125), .Q(n3503)
         );
  OAI22X1 U4168 ( .IN1(n6434), .IN2(n5468), .IN3(n5462), .IN4(n3504), .QN(
        N10376) );
  OA22X1 U4169 ( .IN1(n6434), .IN2(n5440), .IN3(n5445), .IN4(n3505), .Q(n3504)
         );
  OA22X1 U4170 ( .IN1(n5430), .IN2(n3506), .IN3(n6280), .IN4(n5425), .Q(n3505)
         );
  OA22X1 U4171 ( .IN1(n6280), .IN2(n5416), .IN3(n5412), .IN4(n6126), .Q(n3506)
         );
  OAI22X1 U4172 ( .IN1(n6435), .IN2(n5466), .IN3(n5462), .IN4(n3507), .QN(
        N10375) );
  OA22X1 U4173 ( .IN1(n6435), .IN2(n5440), .IN3(n5446), .IN4(n3508), .Q(n3507)
         );
  OA22X1 U4174 ( .IN1(n5430), .IN2(n3509), .IN3(n6281), .IN4(n5425), .Q(n3508)
         );
  OA22X1 U4175 ( .IN1(n6281), .IN2(n5417), .IN3(n5412), .IN4(n6127), .Q(n3509)
         );
  OAI22X1 U4176 ( .IN1(n6436), .IN2(n5467), .IN3(n5462), .IN4(n3510), .QN(
        N10374) );
  OA22X1 U4177 ( .IN1(n6436), .IN2(n5440), .IN3(n5445), .IN4(n3511), .Q(n3510)
         );
  OA22X1 U4178 ( .IN1(n5429), .IN2(n3512), .IN3(n6282), .IN4(n5425), .Q(n3511)
         );
  OA22X1 U4179 ( .IN1(n6282), .IN2(n5418), .IN3(n5412), .IN4(n6128), .Q(n3512)
         );
  OAI22X1 U4180 ( .IN1(n6437), .IN2(n5468), .IN3(n5462), .IN4(n3513), .QN(
        N10373) );
  OA22X1 U4181 ( .IN1(n6437), .IN2(n5439), .IN3(n5445), .IN4(n3514), .Q(n3513)
         );
  OA22X1 U4182 ( .IN1(n5429), .IN2(n3515), .IN3(n6283), .IN4(n5425), .Q(n3514)
         );
  OA22X1 U4183 ( .IN1(n6283), .IN2(n5415), .IN3(n5412), .IN4(n6129), .Q(n3515)
         );
  OAI22X1 U4184 ( .IN1(n6438), .IN2(n5457), .IN3(n5462), .IN4(n3516), .QN(
        N10372) );
  OA22X1 U4185 ( .IN1(n6438), .IN2(n5439), .IN3(n5445), .IN4(n3517), .Q(n3516)
         );
  OA22X1 U4186 ( .IN1(n5429), .IN2(n3518), .IN3(n6284), .IN4(n5425), .Q(n3517)
         );
  OA22X1 U4187 ( .IN1(n6284), .IN2(n5415), .IN3(n5412), .IN4(n6130), .Q(n3518)
         );
  OAI22X1 U4188 ( .IN1(n6439), .IN2(n5456), .IN3(n5462), .IN4(n3519), .QN(
        N10371) );
  OA22X1 U4189 ( .IN1(n6439), .IN2(n5439), .IN3(n5445), .IN4(n3520), .Q(n3519)
         );
  OA22X1 U4190 ( .IN1(n5429), .IN2(n3521), .IN3(n6285), .IN4(n5425), .Q(n3520)
         );
  OA22X1 U4191 ( .IN1(n6285), .IN2(n5421), .IN3(n5412), .IN4(n6131), .Q(n3521)
         );
  OAI22X1 U4192 ( .IN1(n6440), .IN2(n5467), .IN3(n5462), .IN4(n3522), .QN(
        N10370) );
  OA22X1 U4193 ( .IN1(n6440), .IN2(n5439), .IN3(n5445), .IN4(n3523), .Q(n3522)
         );
  OA22X1 U4194 ( .IN1(n5429), .IN2(n3524), .IN3(n6286), .IN4(n5425), .Q(n3523)
         );
  OA22X1 U4195 ( .IN1(n6286), .IN2(n5414), .IN3(n5412), .IN4(n6132), .Q(n3524)
         );
  OAI22X1 U4196 ( .IN1(n6441), .IN2(n5463), .IN3(n5462), .IN4(n3525), .QN(
        N10369) );
  OA22X1 U4197 ( .IN1(n6441), .IN2(n5439), .IN3(n5446), .IN4(n3526), .Q(n3525)
         );
  OA22X1 U4198 ( .IN1(n5429), .IN2(n3527), .IN3(n6287), .IN4(n5425), .Q(n3526)
         );
  OA22X1 U4199 ( .IN1(n6287), .IN2(n5418), .IN3(n5412), .IN4(n6133), .Q(n3527)
         );
  OAI22X1 U4200 ( .IN1(n6442), .IN2(n5463), .IN3(n5462), .IN4(n3528), .QN(
        N10368) );
  OA22X1 U4201 ( .IN1(n6442), .IN2(n5439), .IN3(n5446), .IN4(n3529), .Q(n3528)
         );
  OA22X1 U4202 ( .IN1(n5429), .IN2(n3530), .IN3(n6288), .IN4(n5425), .Q(n3529)
         );
  OA22X1 U4203 ( .IN1(n6288), .IN2(n5417), .IN3(n5271), .IN4(n6134), .Q(n3530)
         );
  OAI22X1 U4204 ( .IN1(n6443), .IN2(n5463), .IN3(n5462), .IN4(n3531), .QN(
        N10366) );
  OA22X1 U4205 ( .IN1(n6443), .IN2(n5439), .IN3(n5446), .IN4(n3532), .Q(n3531)
         );
  OA22X1 U4206 ( .IN1(n5429), .IN2(n3533), .IN3(n6289), .IN4(n5425), .Q(n3532)
         );
  OA22X1 U4207 ( .IN1(n6289), .IN2(n5419), .IN3(n5271), .IN4(n6135), .Q(n3533)
         );
  OAI22X1 U4208 ( .IN1(n6444), .IN2(n5463), .IN3(n5462), .IN4(n3534), .QN(
        N10365) );
  OA22X1 U4209 ( .IN1(n6444), .IN2(n5439), .IN3(n5446), .IN4(n3535), .Q(n3534)
         );
  OA22X1 U4210 ( .IN1(n5429), .IN2(n3536), .IN3(n6290), .IN4(n5425), .Q(n3535)
         );
  OA22X1 U4211 ( .IN1(n6290), .IN2(n5421), .IN3(n5271), .IN4(n6136), .Q(n3536)
         );
  OAI22X1 U4212 ( .IN1(n6445), .IN2(n5463), .IN3(n5462), .IN4(n3537), .QN(
        N10364) );
  OA22X1 U4213 ( .IN1(n6445), .IN2(n5439), .IN3(n5446), .IN4(n3538), .Q(n3537)
         );
  OA22X1 U4214 ( .IN1(n5429), .IN2(n3539), .IN3(n6291), .IN4(n5425), .Q(n3538)
         );
  OA22X1 U4215 ( .IN1(n6291), .IN2(n5418), .IN3(n5271), .IN4(n6137), .Q(n3539)
         );
  OAI22X1 U4216 ( .IN1(n6446), .IN2(n5463), .IN3(n5462), .IN4(n3540), .QN(
        N10363) );
  OA22X1 U4217 ( .IN1(n6446), .IN2(n5439), .IN3(n5447), .IN4(n3541), .Q(n3540)
         );
  OA22X1 U4218 ( .IN1(n5429), .IN2(n3542), .IN3(n6292), .IN4(n5425), .Q(n3541)
         );
  OA22X1 U4219 ( .IN1(n6292), .IN2(n5419), .IN3(n5271), .IN4(n6138), .Q(n3542)
         );
  OAI22X1 U4220 ( .IN1(n6447), .IN2(n5463), .IN3(n5462), .IN4(n3543), .QN(
        N10362) );
  OA22X1 U4221 ( .IN1(n6447), .IN2(n5439), .IN3(n5447), .IN4(n3544), .Q(n3543)
         );
  OA22X1 U4222 ( .IN1(n5429), .IN2(n3545), .IN3(n6293), .IN4(n5425), .Q(n3544)
         );
  OA22X1 U4223 ( .IN1(n6293), .IN2(n5414), .IN3(n5271), .IN4(n6139), .Q(n3545)
         );
  OAI22X1 U4224 ( .IN1(n6448), .IN2(n5467), .IN3(n5462), .IN4(n3546), .QN(
        N10361) );
  OA22X1 U4225 ( .IN1(n6448), .IN2(n5439), .IN3(n5447), .IN4(n3547), .Q(n3546)
         );
  OA22X1 U4226 ( .IN1(n5428), .IN2(n3548), .IN3(n6294), .IN4(n5425), .Q(n3547)
         );
  OA22X1 U4227 ( .IN1(n6294), .IN2(n5414), .IN3(n5271), .IN4(n6140), .Q(n3548)
         );
  OAI22X1 U4228 ( .IN1(n6449), .IN2(n5456), .IN3(n5462), .IN4(n3549), .QN(
        N10360) );
  OA22X1 U4229 ( .IN1(n6449), .IN2(n5439), .IN3(n5447), .IN4(n3550), .Q(n3549)
         );
  OA22X1 U4230 ( .IN1(n5428), .IN2(n3551), .IN3(n6295), .IN4(n5425), .Q(n3550)
         );
  OA22X1 U4231 ( .IN1(n6295), .IN2(n5421), .IN3(n5271), .IN4(n6141), .Q(n3551)
         );
  OAI22X1 U4232 ( .IN1(n6450), .IN2(n5463), .IN3(n5462), .IN4(n3552), .QN(
        N10359) );
  OA22X1 U4233 ( .IN1(n6450), .IN2(n5439), .IN3(n5447), .IN4(n3553), .Q(n3552)
         );
  OA22X1 U4234 ( .IN1(n5428), .IN2(n3554), .IN3(n6296), .IN4(n5425), .Q(n3553)
         );
  OA22X1 U4235 ( .IN1(n6296), .IN2(n5420), .IN3(n5271), .IN4(n6142), .Q(n3554)
         );
  OAI22X1 U4236 ( .IN1(n6451), .IN2(n5457), .IN3(n5462), .IN4(n3555), .QN(
        N10358) );
  OA22X1 U4237 ( .IN1(n6451), .IN2(n5438), .IN3(n5448), .IN4(n3556), .Q(n3555)
         );
  OA22X1 U4238 ( .IN1(n5428), .IN2(n3557), .IN3(n6297), .IN4(n5425), .Q(n3556)
         );
  OA22X1 U4239 ( .IN1(n6297), .IN2(n5420), .IN3(n5271), .IN4(n6143), .Q(n3557)
         );
  OAI22X1 U4240 ( .IN1(n6452), .IN2(n5468), .IN3(n5462), .IN4(n3558), .QN(
        N10357) );
  OA22X1 U4241 ( .IN1(n6452), .IN2(n5438), .IN3(n5448), .IN4(n3559), .Q(n3558)
         );
  OA22X1 U4242 ( .IN1(n5428), .IN2(n3560), .IN3(n6298), .IN4(n5425), .Q(n3559)
         );
  OA22X1 U4243 ( .IN1(n6298), .IN2(n5418), .IN3(n5271), .IN4(n6144), .Q(n3560)
         );
  OAI22X1 U4244 ( .IN1(n6453), .IN2(n5464), .IN3(n5462), .IN4(n3561), .QN(
        N10356) );
  OA22X1 U4245 ( .IN1(n6453), .IN2(n5438), .IN3(n5448), .IN4(n3562), .Q(n3561)
         );
  OA22X1 U4246 ( .IN1(n5428), .IN2(n3563), .IN3(n6299), .IN4(n5425), .Q(n3562)
         );
  OA22X1 U4247 ( .IN1(n6299), .IN2(n5419), .IN3(n5271), .IN4(n6145), .Q(n3563)
         );
  OAI22X1 U4248 ( .IN1(n6454), .IN2(n5466), .IN3(n5459), .IN4(n3564), .QN(
        N10355) );
  OA22X1 U4249 ( .IN1(n6454), .IN2(n5438), .IN3(n5448), .IN4(n3565), .Q(n3564)
         );
  OA22X1 U4250 ( .IN1(n5428), .IN2(n3566), .IN3(n6300), .IN4(n5425), .Q(n3565)
         );
  OA22X1 U4251 ( .IN1(n6300), .IN2(n5420), .IN3(n5271), .IN4(n6146), .Q(n3566)
         );
  OA22X1 U4253 ( .IN1(n6320), .IN2(n5438), .IN3(n5448), .IN4(n3568), .Q(n3567)
         );
  OA22X1 U4257 ( .IN1(n6321), .IN2(n5438), .IN3(n5449), .IN4(n3571), .Q(n3570)
         );
  OA22X1 U4261 ( .IN1(n6322), .IN2(n5438), .IN3(n5449), .IN4(n3574), .Q(n3573)
         );
  OA22X1 U4265 ( .IN1(n6323), .IN2(n5438), .IN3(n5449), .IN4(n3577), .Q(n3576)
         );
  OA22X1 U4269 ( .IN1(n6324), .IN2(n5438), .IN3(n5449), .IN4(n3580), .Q(n3579)
         );
  OA22X1 U4273 ( .IN1(n6325), .IN2(n5438), .IN3(n5449), .IN4(n3583), .Q(n3582)
         );
  OA22X1 U4277 ( .IN1(n6326), .IN2(n5438), .IN3(n5450), .IN4(n3586), .Q(n3585)
         );
  OA22X1 U4281 ( .IN1(n6327), .IN2(n5438), .IN3(n5450), .IN4(n3589), .Q(n3588)
         );
  OA22X1 U4285 ( .IN1(n6328), .IN2(n5438), .IN3(n5450), .IN4(n3592), .Q(n3591)
         );
  OA22X1 U4289 ( .IN1(n6329), .IN2(n5438), .IN3(n5450), .IN4(n3595), .Q(n3594)
         );
  OA22X1 U4293 ( .IN1(n6330), .IN2(n5437), .IN3(n5450), .IN4(n3598), .Q(n3597)
         );
  OA22X1 U4297 ( .IN1(n6331), .IN2(n5437), .IN3(n5451), .IN4(n3601), .Q(n3600)
         );
  OA22X1 U4301 ( .IN1(n6332), .IN2(n5437), .IN3(n5451), .IN4(n3604), .Q(n3603)
         );
  OA22X1 U4305 ( .IN1(n6333), .IN2(n5437), .IN3(n5451), .IN4(n3607), .Q(n3606)
         );
  OA22X1 U4309 ( .IN1(n6334), .IN2(n5437), .IN3(n5451), .IN4(n3610), .Q(n3609)
         );
  OA22X1 U4313 ( .IN1(n6335), .IN2(n5437), .IN3(n5451), .IN4(n3613), .Q(n3612)
         );
  OA22X1 U4317 ( .IN1(n6336), .IN2(n5437), .IN3(n5452), .IN4(n3616), .Q(n3615)
         );
  OA22X1 U4321 ( .IN1(n6337), .IN2(n5437), .IN3(n5452), .IN4(n3619), .Q(n3618)
         );
  OA22X1 U4325 ( .IN1(n6338), .IN2(n5437), .IN3(n5452), .IN4(n3622), .Q(n3621)
         );
  OA22X1 U4329 ( .IN1(n6339), .IN2(n5437), .IN3(n5452), .IN4(n3625), .Q(n3624)
         );
  OA22X1 U4333 ( .IN1(n6340), .IN2(n5437), .IN3(n5452), .IN4(n3628), .Q(n3627)
         );
  OA22X1 U4337 ( .IN1(n6341), .IN2(n5437), .IN3(n5448), .IN4(n3631), .Q(n3630)
         );
  OA22X1 U4341 ( .IN1(n6342), .IN2(n5437), .IN3(n5453), .IN4(n3634), .Q(n3633)
         );
  OA22X1 U4345 ( .IN1(n6343), .IN2(n5437), .IN3(n5454), .IN4(n3637), .Q(n3636)
         );
  OA22X1 U4349 ( .IN1(n6344), .IN2(n5436), .IN3(n5450), .IN4(n3640), .Q(n3639)
         );
  OA22X1 U4353 ( .IN1(n6345), .IN2(n5436), .IN3(n5447), .IN4(n3643), .Q(n3642)
         );
  OA22X1 U4357 ( .IN1(n6346), .IN2(n5436), .IN3(n5449), .IN4(n3646), .Q(n3645)
         );
  OA22X1 U4361 ( .IN1(n6315), .IN2(n5436), .IN3(n5450), .IN4(n3649), .Q(n3648)
         );
  OA22X1 U4365 ( .IN1(n6316), .IN2(n5436), .IN3(n5445), .IN4(n3652), .Q(n3651)
         );
  OA22X1 U4369 ( .IN1(n6317), .IN2(n5436), .IN3(n5446), .IN4(n3655), .Q(n3654)
         );
  OA22X1 U4373 ( .IN1(n6318), .IN2(n5436), .IN3(n5447), .IN4(n3658), .Q(n3657)
         );
  OA22X1 U4377 ( .IN1(n6319), .IN2(n5436), .IN3(n5452), .IN4(n3661), .Q(n3660)
         );
  OAI22X1 U4380 ( .IN1(n6455), .IN2(n5465), .IN3(n5458), .IN4(n3663), .QN(
        N10322) );
  OA22X1 U4381 ( .IN1(n6455), .IN2(n5436), .IN3(n5451), .IN4(n3664), .Q(n3663)
         );
  OA22X1 U4382 ( .IN1(n5428), .IN2(n3665), .IN3(n6301), .IN4(n5424), .Q(n3664)
         );
  OA22X1 U4383 ( .IN1(n6301), .IN2(n5415), .IN3(n5271), .IN4(n6147), .Q(n3665)
         );
  OAI22X1 U4384 ( .IN1(n6456), .IN2(n5464), .IN3(n5459), .IN4(n3666), .QN(
        N10321) );
  OA22X1 U4385 ( .IN1(n6456), .IN2(n5436), .IN3(n5449), .IN4(n3667), .Q(n3666)
         );
  OA22X1 U4386 ( .IN1(n5428), .IN2(n3668), .IN3(n6302), .IN4(n5424), .Q(n3667)
         );
  OA22X1 U4387 ( .IN1(n6302), .IN2(n5421), .IN3(n5271), .IN4(n6148), .Q(n3668)
         );
  OAI22X1 U4388 ( .IN1(n6457), .IN2(n5457), .IN3(n5458), .IN4(n3669), .QN(
        N10320) );
  OA22X1 U4389 ( .IN1(n6457), .IN2(n5436), .IN3(n5449), .IN4(n3670), .Q(n3669)
         );
  OA22X1 U4390 ( .IN1(n5428), .IN2(n3671), .IN3(n6303), .IN4(n5424), .Q(n3670)
         );
  OA22X1 U4391 ( .IN1(n6303), .IN2(n5416), .IN3(n5271), .IN4(n6149), .Q(n3671)
         );
  OAI22X1 U4392 ( .IN1(n6458), .IN2(n5468), .IN3(n5459), .IN4(n3672), .QN(
        N10319) );
  OA22X1 U4393 ( .IN1(n6458), .IN2(n5436), .IN3(n5453), .IN4(n3673), .Q(n3672)
         );
  OA22X1 U4394 ( .IN1(n5428), .IN2(n3674), .IN3(n6304), .IN4(n5424), .Q(n3673)
         );
  OA22X1 U4395 ( .IN1(n6304), .IN2(n5420), .IN3(n5271), .IN4(n6150), .Q(n3674)
         );
  OAI22X1 U4396 ( .IN1(n6459), .IN2(n5465), .IN3(n5458), .IN4(n3675), .QN(
        N10318) );
  OA22X1 U4397 ( .IN1(n6459), .IN2(n5436), .IN3(n5453), .IN4(n3676), .Q(n3675)
         );
  OA22X1 U4398 ( .IN1(n5428), .IN2(n3677), .IN3(n6305), .IN4(n5424), .Q(n3676)
         );
  OA22X1 U4399 ( .IN1(n6305), .IN2(n5416), .IN3(n5412), .IN4(n6151), .Q(n3677)
         );
  NAND4X0 U4400 ( .IN1(n3678), .IN2(n5436), .IN3(n3679), .IN4(n5424), .QN(
        decodedVector_o[5]) );
  NAND4X0 U4402 ( .IN1(decodedPacketValid[4]), .IN2(N2172), .IN3(n2908), .IN4(
        n5990), .QN(n3302) );
  NAND4X0 U4403 ( .IN1(decodedPacketValid[7]), .IN2(N8580), .IN3(n2909), .IN4(
        n5987), .QN(n3296) );
  NAND4X0 U4404 ( .IN1(decodedPacketValid[6]), .IN2(N6444), .IN3(n2910), .IN4(
        n5988), .QN(n3298) );
  NAND4X0 U4405 ( .IN1(decodedPacketValid[3]), .IN2(N1068), .IN3(N1070), .IN4(
        n5991), .QN(n3678) );
  OA22X1 U4423 ( .IN1(n5856), .IN2(n5385), .IN3(n5389), .IN4(n3697), .Q(n3696)
         );
  OAI22X1 U4426 ( .IN1(n6384), .IN2(n5409), .IN3(n5401), .IN4(n3699), .QN(
        N10311) );
  OA22X1 U4427 ( .IN1(n6349), .IN2(n5385), .IN3(n5395), .IN4(n3700), .Q(n3699)
         );
  OA22X1 U4428 ( .IN1(n5376), .IN2(n3701), .IN3(n6230), .IN4(n5368), .Q(n3700)
         );
  OA22X1 U4429 ( .IN1(n6195), .IN2(n5355), .IN3(n5269), .IN4(n6076), .Q(n3701)
         );
  OAI22X1 U4430 ( .IN1(n6376), .IN2(n5409), .IN3(n5401), .IN4(n3702), .QN(
        N10310) );
  OA22X1 U4431 ( .IN1(n6348), .IN2(n5385), .IN3(n5389), .IN4(n3703), .Q(n3702)
         );
  OA22X1 U4432 ( .IN1(n5376), .IN2(n3704), .IN3(n6222), .IN4(n5368), .Q(n3703)
         );
  OA22X1 U4433 ( .IN1(n6194), .IN2(n5355), .IN3(n5354), .IN4(n6068), .Q(n3704)
         );
  OAI22X1 U4434 ( .IN1(n6372), .IN2(n5409), .IN3(n5401), .IN4(n3705), .QN(
        N10309) );
  OA22X1 U4435 ( .IN1(n6374), .IN2(n5385), .IN3(n5386), .IN4(n3706), .Q(n3705)
         );
  OA22X1 U4436 ( .IN1(n5376), .IN2(n3707), .IN3(n6218), .IN4(n5368), .Q(n3706)
         );
  OA22X1 U4437 ( .IN1(n6220), .IN2(n5355), .IN3(n5354), .IN4(n6065), .Q(n3707)
         );
  OA22X1 U4439 ( .IN1(n6371), .IN2(n5385), .IN3(n5393), .IN4(n3709), .Q(n3708)
         );
  OAI22X1 U4442 ( .IN1(n6373), .IN2(n5409), .IN3(n5401), .IN4(n3711), .QN(
        N10307) );
  OA22X1 U4443 ( .IN1(n6370), .IN2(n5385), .IN3(n5392), .IN4(n3712), .Q(n3711)
         );
  OA22X1 U4444 ( .IN1(n5376), .IN2(n3713), .IN3(n6219), .IN4(n5368), .Q(n3712)
         );
  OA22X1 U4445 ( .IN1(n6216), .IN2(n5355), .IN3(n5354), .IN4(n6065), .Q(n3713)
         );
  OAI22X1 U4446 ( .IN1(n6395), .IN2(n5409), .IN3(n5402), .IN4(n3714), .QN(
        N10306) );
  OA22X1 U4447 ( .IN1(n6347), .IN2(n5385), .IN3(n5391), .IN4(n3715), .Q(n3714)
         );
  OA22X1 U4448 ( .IN1(n5375), .IN2(n3716), .IN3(n6245), .IN4(n5368), .Q(n3715)
         );
  OA22X1 U4449 ( .IN1(n6193), .IN2(n5355), .IN3(n5354), .IN4(n6091), .Q(n3716)
         );
  OAI22X1 U4450 ( .IN1(n5967), .IN2(n5409), .IN3(n5402), .IN4(n3717), .QN(
        N10305) );
  OA22X1 U4451 ( .IN1(n6369), .IN2(n5385), .IN3(n5386), .IN4(n3718), .Q(n3717)
         );
  OA22X1 U4452 ( .IN1(n5375), .IN2(n3719), .IN3(n5952), .IN4(n5368), .Q(n3718)
         );
  OA22X1 U4453 ( .IN1(n6215), .IN2(n5356), .IN3(n5354), .IN4(n5937), .Q(n3719)
         );
  OAI22X1 U4454 ( .IN1(n5968), .IN2(n5408), .IN3(n5402), .IN4(n3720), .QN(
        N10304) );
  OA22X1 U4455 ( .IN1(n6368), .IN2(n5385), .IN3(n5387), .IN4(n3721), .Q(n3720)
         );
  OA22X1 U4456 ( .IN1(n5375), .IN2(n3722), .IN3(n5953), .IN4(n5368), .Q(n3721)
         );
  OA22X1 U4457 ( .IN1(n6214), .IN2(n5356), .IN3(n5354), .IN4(n5938), .Q(n3722)
         );
  OAI22X1 U4458 ( .IN1(n5969), .IN2(n5408), .IN3(n5402), .IN4(n3723), .QN(
        N10303) );
  OA22X1 U4459 ( .IN1(n6367), .IN2(n5385), .IN3(n5388), .IN4(n3724), .Q(n3723)
         );
  OA22X1 U4460 ( .IN1(n5375), .IN2(n3725), .IN3(n5954), .IN4(n5368), .Q(n3724)
         );
  OA22X1 U4461 ( .IN1(n6213), .IN2(n5356), .IN3(n5354), .IN4(n5939), .Q(n3725)
         );
  OAI22X1 U4462 ( .IN1(n5970), .IN2(n5408), .IN3(n5402), .IN4(n3726), .QN(
        N10302) );
  OA22X1 U4463 ( .IN1(n6366), .IN2(n5385), .IN3(n5396), .IN4(n3727), .Q(n3726)
         );
  OA22X1 U4464 ( .IN1(n5375), .IN2(n3728), .IN3(n5955), .IN4(n5368), .Q(n3727)
         );
  OA22X1 U4465 ( .IN1(n6212), .IN2(n5356), .IN3(n5354), .IN4(n5940), .Q(n3728)
         );
  OAI22X1 U4466 ( .IN1(n5971), .IN2(n5408), .IN3(n5402), .IN4(n3729), .QN(
        N10301) );
  OA22X1 U4467 ( .IN1(n6365), .IN2(n5384), .IN3(n5390), .IN4(n3730), .Q(n3729)
         );
  OA22X1 U4468 ( .IN1(n5375), .IN2(n3731), .IN3(n5956), .IN4(n5368), .Q(n3730)
         );
  OA22X1 U4469 ( .IN1(n6211), .IN2(n5356), .IN3(n5354), .IN4(n5941), .Q(n3731)
         );
  OAI22X1 U4470 ( .IN1(n5972), .IN2(n5408), .IN3(n5402), .IN4(n3732), .QN(
        N10300) );
  OA22X1 U4471 ( .IN1(n6364), .IN2(n5384), .IN3(n5393), .IN4(n3733), .Q(n3732)
         );
  OA22X1 U4472 ( .IN1(n5375), .IN2(n3734), .IN3(n5957), .IN4(n5368), .Q(n3733)
         );
  OA22X1 U4473 ( .IN1(n6210), .IN2(n5357), .IN3(n5354), .IN4(n5942), .Q(n3734)
         );
  OAI22X1 U4474 ( .IN1(n5973), .IN2(n5408), .IN3(n5402), .IN4(n3735), .QN(
        N10299) );
  OA22X1 U4475 ( .IN1(n6363), .IN2(n5384), .IN3(n5392), .IN4(n3736), .Q(n3735)
         );
  OA22X1 U4476 ( .IN1(n5375), .IN2(n3737), .IN3(n5958), .IN4(n5368), .Q(n3736)
         );
  OA22X1 U4477 ( .IN1(n6209), .IN2(n5357), .IN3(n5354), .IN4(n5943), .Q(n3737)
         );
  OAI22X1 U4478 ( .IN1(n5974), .IN2(n5408), .IN3(n5402), .IN4(n3738), .QN(
        N10298) );
  OA22X1 U4479 ( .IN1(n6362), .IN2(n5384), .IN3(n5396), .IN4(n3739), .Q(n3738)
         );
  OA22X1 U4480 ( .IN1(n5375), .IN2(n3740), .IN3(n5959), .IN4(n5368), .Q(n3739)
         );
  OA22X1 U4481 ( .IN1(n6208), .IN2(n5357), .IN3(n5354), .IN4(n5944), .Q(n3740)
         );
  OAI22X1 U4482 ( .IN1(n5975), .IN2(n5405), .IN3(n5402), .IN4(n3741), .QN(
        N10297) );
  OA22X1 U4483 ( .IN1(n6308), .IN2(n5384), .IN3(n5395), .IN4(n3742), .Q(n3741)
         );
  OA22X1 U4484 ( .IN1(n5375), .IN2(n3743), .IN3(n5960), .IN4(n5367), .Q(n3742)
         );
  OA22X1 U4485 ( .IN1(n6154), .IN2(n5357), .IN3(n5354), .IN4(n5945), .Q(n3743)
         );
  OAI22X1 U4486 ( .IN1(n5976), .IN2(n5408), .IN3(n5402), .IN4(n3744), .QN(
        N10296) );
  OA22X1 U4487 ( .IN1(n6309), .IN2(n5384), .IN3(n5386), .IN4(n3745), .Q(n3744)
         );
  OA22X1 U4488 ( .IN1(n5375), .IN2(n3746), .IN3(n5961), .IN4(n5367), .Q(n3745)
         );
  OA22X1 U4489 ( .IN1(n6155), .IN2(n5357), .IN3(n5354), .IN4(n5946), .Q(n3746)
         );
  OAI22X1 U4490 ( .IN1(n5977), .IN2(n5398), .IN3(n5402), .IN4(n3747), .QN(
        N10295) );
  OA22X1 U4491 ( .IN1(n6310), .IN2(n5384), .IN3(n5389), .IN4(n3748), .Q(n3747)
         );
  OA22X1 U4492 ( .IN1(n5375), .IN2(n3749), .IN3(n5962), .IN4(n5367), .Q(n3748)
         );
  OA22X1 U4493 ( .IN1(n6156), .IN2(n5358), .IN3(n5354), .IN4(n5947), .Q(n3749)
         );
  OAI22X1 U4494 ( .IN1(n5978), .IN2(n5405), .IN3(n5402), .IN4(n3750), .QN(
        N10294) );
  OA22X1 U4495 ( .IN1(n6311), .IN2(n5384), .IN3(n5396), .IN4(n3751), .Q(n3750)
         );
  OA22X1 U4496 ( .IN1(n5374), .IN2(n3752), .IN3(n5963), .IN4(n5367), .Q(n3751)
         );
  OA22X1 U4497 ( .IN1(n6157), .IN2(n5358), .IN3(n5354), .IN4(n5948), .Q(n3752)
         );
  OAI22X1 U4498 ( .IN1(n5979), .IN2(n5404), .IN3(n5402), .IN4(n3753), .QN(
        N10293) );
  OA22X1 U4499 ( .IN1(n6312), .IN2(n5384), .IN3(n5395), .IN4(n3754), .Q(n3753)
         );
  OA22X1 U4500 ( .IN1(n5374), .IN2(n3755), .IN3(n5964), .IN4(n5367), .Q(n3754)
         );
  OA22X1 U4501 ( .IN1(n6158), .IN2(n5358), .IN3(n5354), .IN4(n5949), .Q(n3755)
         );
  OAI22X1 U4502 ( .IN1(n5980), .IN2(n5407), .IN3(n5402), .IN4(n3756), .QN(
        N10292) );
  OA22X1 U4503 ( .IN1(n6313), .IN2(n5384), .IN3(n5394), .IN4(n3757), .Q(n3756)
         );
  OA22X1 U4504 ( .IN1(n5374), .IN2(n3758), .IN3(n5965), .IN4(n5367), .Q(n3757)
         );
  OA22X1 U4505 ( .IN1(n6159), .IN2(n5358), .IN3(n5354), .IN4(n5950), .Q(n3758)
         );
  OAI22X1 U4506 ( .IN1(n5981), .IN2(n5409), .IN3(n5402), .IN4(n3759), .QN(
        N10291) );
  OA22X1 U4507 ( .IN1(n6314), .IN2(n5384), .IN3(n5395), .IN4(n3760), .Q(n3759)
         );
  OA22X1 U4508 ( .IN1(n5374), .IN2(n3761), .IN3(n5966), .IN4(n5367), .Q(n3760)
         );
  OA22X1 U4509 ( .IN1(n6160), .IN2(n5358), .IN3(n5354), .IN4(n5951), .Q(n3761)
         );
  OAI22X1 U4510 ( .IN1(n6375), .IN2(n5408), .IN3(n5402), .IN4(n3762), .QN(
        N10290) );
  OA22X1 U4511 ( .IN1(n6307), .IN2(n5384), .IN3(n5394), .IN4(n3763), .Q(n3762)
         );
  OA22X1 U4512 ( .IN1(n5374), .IN2(n3764), .IN3(n6221), .IN4(n5367), .Q(n3763)
         );
  OA22X1 U4513 ( .IN1(n6153), .IN2(n5359), .IN3(n5354), .IN4(n6067), .Q(n3764)
         );
  OAI22X1 U4514 ( .IN1(n6372), .IN2(n5406), .IN3(n5402), .IN4(n3765), .QN(
        N10288) );
  OA22X1 U4515 ( .IN1(n6306), .IN2(n5384), .IN3(n5395), .IN4(n3766), .Q(n3765)
         );
  OA22X1 U4516 ( .IN1(n5374), .IN2(n3767), .IN3(n6218), .IN4(n5367), .Q(n3766)
         );
  OA22X1 U4517 ( .IN1(n6152), .IN2(n5359), .IN3(n5354), .IN4(n6064), .Q(n3767)
         );
  OAI22X1 U4518 ( .IN1(n6377), .IN2(n5398), .IN3(n5402), .IN4(n3768), .QN(
        N10286) );
  OA22X1 U4519 ( .IN1(n6422), .IN2(n5384), .IN3(n5396), .IN4(n3769), .Q(n3768)
         );
  OA22X1 U4520 ( .IN1(n5374), .IN2(n3770), .IN3(n6223), .IN4(n5367), .Q(n3769)
         );
  OA22X1 U4521 ( .IN1(n6268), .IN2(n5359), .IN3(n5354), .IN4(n6069), .Q(n3770)
         );
  OAI22X1 U4522 ( .IN1(n6378), .IN2(n5404), .IN3(n5402), .IN4(n3771), .QN(
        N10285) );
  OA22X1 U4523 ( .IN1(n6421), .IN2(n5383), .IN3(n5392), .IN4(n3772), .Q(n3771)
         );
  OA22X1 U4524 ( .IN1(n5374), .IN2(n3773), .IN3(n6224), .IN4(n5367), .Q(n3772)
         );
  OA22X1 U4525 ( .IN1(n6267), .IN2(n5359), .IN3(n5354), .IN4(n6070), .Q(n3773)
         );
  OAI22X1 U4526 ( .IN1(n6379), .IN2(n5407), .IN3(n5402), .IN4(n3774), .QN(
        N10284) );
  OA22X1 U4527 ( .IN1(n6420), .IN2(n5383), .IN3(n5389), .IN4(n3775), .Q(n3774)
         );
  OA22X1 U4528 ( .IN1(n5374), .IN2(n3776), .IN3(n6225), .IN4(n5367), .Q(n3775)
         );
  OA22X1 U4529 ( .IN1(n6266), .IN2(n5359), .IN3(n5354), .IN4(n6071), .Q(n3776)
         );
  OAI22X1 U4530 ( .IN1(n6380), .IN2(n5397), .IN3(n5402), .IN4(n3777), .QN(
        N10283) );
  OA22X1 U4531 ( .IN1(n6419), .IN2(n5383), .IN3(n5394), .IN4(n3778), .Q(n3777)
         );
  OA22X1 U4532 ( .IN1(n5374), .IN2(n3779), .IN3(n6226), .IN4(n5367), .Q(n3778)
         );
  OA22X1 U4533 ( .IN1(n6265), .IN2(n5360), .IN3(n5354), .IN4(n6072), .Q(n3779)
         );
  OAI22X1 U4534 ( .IN1(n6381), .IN2(n5409), .IN3(n5402), .IN4(n3780), .QN(
        N10282) );
  OA22X1 U4535 ( .IN1(n6418), .IN2(n5383), .IN3(n5394), .IN4(n3781), .Q(n3780)
         );
  OA22X1 U4536 ( .IN1(n5374), .IN2(n3782), .IN3(n6227), .IN4(n5367), .Q(n3781)
         );
  OA22X1 U4537 ( .IN1(n6264), .IN2(n5360), .IN3(n5354), .IN4(n6073), .Q(n3782)
         );
  OAI22X1 U4538 ( .IN1(n6382), .IN2(n5407), .IN3(n5402), .IN4(n3783), .QN(
        N10281) );
  OA22X1 U4539 ( .IN1(n6417), .IN2(n5383), .IN3(n5395), .IN4(n3784), .Q(n3783)
         );
  OA22X1 U4540 ( .IN1(n5374), .IN2(n3785), .IN3(n6228), .IN4(n5367), .Q(n3784)
         );
  OA22X1 U4541 ( .IN1(n6263), .IN2(n5360), .IN3(n5354), .IN4(n6074), .Q(n3785)
         );
  OAI22X1 U4542 ( .IN1(n6383), .IN2(n5407), .IN3(n5402), .IN4(n3786), .QN(
        N10280) );
  OA22X1 U4543 ( .IN1(n6416), .IN2(n5383), .IN3(n5396), .IN4(n3787), .Q(n3786)
         );
  OA22X1 U4544 ( .IN1(n5373), .IN2(n3788), .IN3(n6229), .IN4(n5367), .Q(n3787)
         );
  OA22X1 U4545 ( .IN1(n6262), .IN2(n5360), .IN3(n5354), .IN4(n6075), .Q(n3788)
         );
  OAI22X1 U4546 ( .IN1(n6385), .IN2(n5407), .IN3(n5402), .IN4(n3789), .QN(
        N10279) );
  OA22X1 U4547 ( .IN1(n6359), .IN2(n5383), .IN3(n5393), .IN4(n3790), .Q(n3789)
         );
  OA22X1 U4548 ( .IN1(n5373), .IN2(n3791), .IN3(n6231), .IN4(n5367), .Q(n3790)
         );
  OA22X1 U4549 ( .IN1(n6205), .IN2(n5360), .IN3(n5354), .IN4(n6077), .Q(n3791)
         );
  OAI22X1 U4550 ( .IN1(n6386), .IN2(n5407), .IN3(n5402), .IN4(n3792), .QN(
        N10278) );
  OA22X1 U4551 ( .IN1(n6358), .IN2(n5383), .IN3(n5387), .IN4(n3793), .Q(n3792)
         );
  OA22X1 U4552 ( .IN1(n5373), .IN2(n3794), .IN3(n6232), .IN4(n5367), .Q(n3793)
         );
  OA22X1 U4553 ( .IN1(n6204), .IN2(n5359), .IN3(n5354), .IN4(n6078), .Q(n3794)
         );
  OAI22X1 U4554 ( .IN1(n6387), .IN2(n5407), .IN3(n5402), .IN4(n3795), .QN(
        N10277) );
  OA22X1 U4555 ( .IN1(n6357), .IN2(n5383), .IN3(n5389), .IN4(n3796), .Q(n3795)
         );
  OA22X1 U4556 ( .IN1(n5373), .IN2(n3797), .IN3(n6233), .IN4(n5367), .Q(n3796)
         );
  OA22X1 U4557 ( .IN1(n6203), .IN2(n5355), .IN3(n5354), .IN4(n6079), .Q(n3797)
         );
  OAI22X1 U4558 ( .IN1(n6388), .IN2(n5407), .IN3(n5402), .IN4(n3798), .QN(
        N10276) );
  OA22X1 U4559 ( .IN1(n6356), .IN2(n5383), .IN3(n5393), .IN4(n3799), .Q(n3798)
         );
  OA22X1 U4560 ( .IN1(n5373), .IN2(n3800), .IN3(n6234), .IN4(n5367), .Q(n3799)
         );
  OA22X1 U4561 ( .IN1(n6202), .IN2(n5360), .IN3(n5354), .IN4(n6080), .Q(n3800)
         );
  OAI22X1 U4562 ( .IN1(n6389), .IN2(n5407), .IN3(n5402), .IN4(n3801), .QN(
        N10275) );
  OA22X1 U4563 ( .IN1(n6355), .IN2(n5383), .IN3(n5392), .IN4(n3802), .Q(n3801)
         );
  OA22X1 U4564 ( .IN1(n5373), .IN2(n3803), .IN3(n6235), .IN4(n5367), .Q(n3802)
         );
  OA22X1 U4565 ( .IN1(n6201), .IN2(n5355), .IN3(n5353), .IN4(n6081), .Q(n3803)
         );
  OAI22X1 U4566 ( .IN1(n6390), .IN2(n5406), .IN3(n5402), .IN4(n3804), .QN(
        N10274) );
  OA22X1 U4567 ( .IN1(n6354), .IN2(n5383), .IN3(n5390), .IN4(n3805), .Q(n3804)
         );
  OA22X1 U4568 ( .IN1(n5373), .IN2(n3806), .IN3(n6236), .IN4(n5367), .Q(n3805)
         );
  OA22X1 U4569 ( .IN1(n6200), .IN2(n5356), .IN3(n5353), .IN4(n6082), .Q(n3806)
         );
  OAI22X1 U4570 ( .IN1(n6391), .IN2(n5406), .IN3(n5402), .IN4(n3807), .QN(
        N10273) );
  OA22X1 U4571 ( .IN1(n6353), .IN2(n5383), .IN3(n5391), .IN4(n3808), .Q(n3807)
         );
  OA22X1 U4572 ( .IN1(n5373), .IN2(n3809), .IN3(n6237), .IN4(n5367), .Q(n3808)
         );
  OA22X1 U4573 ( .IN1(n6199), .IN2(n5356), .IN3(n5353), .IN4(n6083), .Q(n3809)
         );
  OAI22X1 U4574 ( .IN1(n6400), .IN2(n5406), .IN3(n5402), .IN4(n3810), .QN(
        N10272) );
  OA22X1 U4575 ( .IN1(n6415), .IN2(n5383), .IN3(n5386), .IN4(n3811), .Q(n3810)
         );
  OA22X1 U4576 ( .IN1(n5373), .IN2(n3812), .IN3(n6246), .IN4(n5367), .Q(n3811)
         );
  OA22X1 U4577 ( .IN1(n6261), .IN2(n5357), .IN3(n5353), .IN4(n6092), .Q(n3812)
         );
  OAI22X1 U4578 ( .IN1(n6406), .IN2(n5406), .IN3(n5402), .IN4(n3813), .QN(
        N10271) );
  OA22X1 U4579 ( .IN1(n6414), .IN2(n5382), .IN3(n5387), .IN4(n3814), .Q(n3813)
         );
  OA22X1 U4580 ( .IN1(n5373), .IN2(n3815), .IN3(n6252), .IN4(n5367), .Q(n3814)
         );
  OA22X1 U4581 ( .IN1(n6260), .IN2(n5358), .IN3(n5353), .IN4(n6098), .Q(n3815)
         );
  OAI22X1 U4582 ( .IN1(n6407), .IN2(n5406), .IN3(n5402), .IN4(n3816), .QN(
        N10270) );
  OA22X1 U4583 ( .IN1(n6413), .IN2(n5382), .IN3(n5388), .IN4(n3817), .Q(n3816)
         );
  OA22X1 U4584 ( .IN1(n5373), .IN2(n3818), .IN3(n6253), .IN4(n5367), .Q(n3817)
         );
  OA22X1 U4585 ( .IN1(n6259), .IN2(n5360), .IN3(n5353), .IN4(n6099), .Q(n3818)
         );
  OAI22X1 U4586 ( .IN1(n6408), .IN2(n5406), .IN3(n5402), .IN4(n3819), .QN(
        N10269) );
  OA22X1 U4587 ( .IN1(n6412), .IN2(n5382), .IN3(n5393), .IN4(n3820), .Q(n3819)
         );
  OA22X1 U4588 ( .IN1(n5373), .IN2(n3821), .IN3(n6254), .IN4(n5367), .Q(n3820)
         );
  OA22X1 U4589 ( .IN1(n6258), .IN2(n5358), .IN3(n5353), .IN4(n6100), .Q(n3821)
         );
  OAI22X1 U4590 ( .IN1(n6409), .IN2(n5406), .IN3(n5402), .IN4(n3822), .QN(
        N10268) );
  OA22X1 U4591 ( .IN1(n6411), .IN2(n5382), .IN3(n5387), .IN4(n3823), .Q(n3822)
         );
  OA22X1 U4592 ( .IN1(n5372), .IN2(n3824), .IN3(n6255), .IN4(n5367), .Q(n3823)
         );
  OA22X1 U4593 ( .IN1(n6257), .IN2(n5361), .IN3(n5353), .IN4(n6101), .Q(n3824)
         );
  OAI22X1 U4594 ( .IN1(n6401), .IN2(n5405), .IN3(n5402), .IN4(n3825), .QN(
        N10267) );
  OA22X1 U4595 ( .IN1(n6410), .IN2(n5382), .IN3(n5389), .IN4(n3826), .Q(n3825)
         );
  OA22X1 U4596 ( .IN1(n5372), .IN2(n3827), .IN3(n6247), .IN4(n5367), .Q(n3826)
         );
  OA22X1 U4597 ( .IN1(n6256), .IN2(n5362), .IN3(n5353), .IN4(n6093), .Q(n3827)
         );
  OAI22X1 U4598 ( .IN1(n6399), .IN2(n5405), .IN3(n5402), .IN4(n3828), .QN(
        N10266) );
  OA22X1 U4599 ( .IN1(n6352), .IN2(n5382), .IN3(n5392), .IN4(n3829), .Q(n3828)
         );
  OA22X1 U4600 ( .IN1(n5372), .IN2(n3830), .IN3(n6244), .IN4(n5367), .Q(n3829)
         );
  OA22X1 U4601 ( .IN1(n6198), .IN2(n5355), .IN3(n5353), .IN4(n6090), .Q(n3830)
         );
  OAI22X1 U4602 ( .IN1(n6398), .IN2(n5405), .IN3(n5403), .IN4(n3831), .QN(
        N10265) );
  OA22X1 U4603 ( .IN1(n6402), .IN2(n5382), .IN3(n5386), .IN4(n3832), .Q(n3831)
         );
  OA22X1 U4604 ( .IN1(n5372), .IN2(n3833), .IN3(n6243), .IN4(n5367), .Q(n3832)
         );
  OA22X1 U4605 ( .IN1(n6248), .IN2(n5356), .IN3(n5353), .IN4(n6089), .Q(n3833)
         );
  OAI22X1 U4606 ( .IN1(n6397), .IN2(n5405), .IN3(n5403), .IN4(n3834), .QN(
        N10264) );
  OA22X1 U4607 ( .IN1(n6403), .IN2(n5382), .IN3(n5388), .IN4(n3835), .Q(n3834)
         );
  OA22X1 U4608 ( .IN1(n5372), .IN2(n3836), .IN3(n6242), .IN4(n5367), .Q(n3835)
         );
  OA22X1 U4609 ( .IN1(n6249), .IN2(n5357), .IN3(n5353), .IN4(n6087), .Q(n3836)
         );
  OAI22X1 U4610 ( .IN1(n6396), .IN2(n5405), .IN3(n5403), .IN4(n3837), .QN(
        N10263) );
  OA22X1 U4611 ( .IN1(n6404), .IN2(n5382), .IN3(n5390), .IN4(n3838), .Q(n3837)
         );
  OA22X1 U4612 ( .IN1(n5372), .IN2(n3839), .IN3(n6241), .IN4(n5367), .Q(n3838)
         );
  OA22X1 U4613 ( .IN1(n6250), .IN2(n5360), .IN3(n5353), .IN4(n6088), .Q(n3839)
         );
  OAI22X1 U4614 ( .IN1(n6398), .IN2(n5405), .IN3(n5403), .IN4(n3840), .QN(
        N10262) );
  OA22X1 U4615 ( .IN1(n6405), .IN2(n5382), .IN3(n5387), .IN4(n3841), .Q(n3840)
         );
  OA22X1 U4616 ( .IN1(n5372), .IN2(n3842), .IN3(n6245), .IN4(n5367), .Q(n3841)
         );
  OA22X1 U4617 ( .IN1(n6251), .IN2(n5361), .IN3(n5353), .IN4(n6087), .Q(n3842)
         );
  OAI22X1 U4618 ( .IN1(n6394), .IN2(n5405), .IN3(n5403), .IN4(n3843), .QN(
        N10261) );
  OA22X1 U4619 ( .IN1(n6393), .IN2(n5382), .IN3(n5396), .IN4(n3844), .Q(n3843)
         );
  OA22X1 U4620 ( .IN1(n5372), .IN2(n3845), .IN3(n6240), .IN4(n5367), .Q(n3844)
         );
  OA22X1 U4621 ( .IN1(n6239), .IN2(n5362), .IN3(n5353), .IN4(n6086), .Q(n3845)
         );
  OAI22X1 U4622 ( .IN1(n6361), .IN2(n5404), .IN3(n5403), .IN4(n3846), .QN(
        N10260) );
  OA22X1 U4623 ( .IN1(n6360), .IN2(n5382), .IN3(n5392), .IN4(n3847), .Q(n3846)
         );
  OA22X1 U4624 ( .IN1(n5372), .IN2(n3848), .IN3(n6207), .IN4(n5366), .Q(n3847)
         );
  OA22X1 U4625 ( .IN1(n6206), .IN2(n5355), .IN3(n5353), .IN4(n6053), .Q(n3848)
         );
  OAI22X1 U4626 ( .IN1(n6350), .IN2(n5404), .IN3(n5403), .IN4(n3849), .QN(
        N10259) );
  OA22X1 U4627 ( .IN1(n6351), .IN2(n5382), .IN3(n5392), .IN4(n3850), .Q(n3849)
         );
  OA22X1 U4628 ( .IN1(n5372), .IN2(n3851), .IN3(n6196), .IN4(n5366), .Q(n3850)
         );
  OA22X1 U4629 ( .IN1(n6197), .IN2(n5356), .IN3(n5353), .IN4(n6042), .Q(n3851)
         );
  OAI22X1 U4630 ( .IN1(n6395), .IN2(n5404), .IN3(n5403), .IN4(n3852), .QN(
        N10258) );
  OA22X1 U4631 ( .IN1(n6392), .IN2(n5382), .IN3(n5393), .IN4(n3853), .Q(n3852)
         );
  OA22X1 U4632 ( .IN1(n5372), .IN2(n3854), .IN3(n6241), .IN4(n5366), .Q(n3853)
         );
  OA22X1 U4633 ( .IN1(n6238), .IN2(n5361), .IN3(n5353), .IN4(n6087), .Q(n3854)
         );
  OAI22X1 U4634 ( .IN1(n6423), .IN2(n5404), .IN3(n5403), .IN4(n3855), .QN(
        N10257) );
  OA22X1 U4635 ( .IN1(n6423), .IN2(n5381), .IN3(n5394), .IN4(n3856), .Q(n3855)
         );
  OA22X1 U4636 ( .IN1(n5372), .IN2(n3857), .IN3(n6269), .IN4(n5366), .Q(n3856)
         );
  OA22X1 U4637 ( .IN1(n6269), .IN2(n5361), .IN3(n5353), .IN4(n6115), .Q(n3857)
         );
  OAI22X1 U4638 ( .IN1(n6424), .IN2(n5404), .IN3(n5403), .IN4(n3858), .QN(
        N10256) );
  OA22X1 U4639 ( .IN1(n6424), .IN2(n5381), .IN3(n5389), .IN4(n3859), .Q(n3858)
         );
  OA22X1 U4640 ( .IN1(n5371), .IN2(n3860), .IN3(n6270), .IN4(n5366), .Q(n3859)
         );
  OA22X1 U4641 ( .IN1(n6270), .IN2(n5361), .IN3(n5353), .IN4(n6116), .Q(n3860)
         );
  OAI22X1 U4642 ( .IN1(n6425), .IN2(n5404), .IN3(n5403), .IN4(n3861), .QN(
        N10255) );
  OA22X1 U4643 ( .IN1(n6425), .IN2(n5381), .IN3(n5394), .IN4(n3862), .Q(n3861)
         );
  OA22X1 U4644 ( .IN1(n5371), .IN2(n3863), .IN3(n6271), .IN4(n5366), .Q(n3862)
         );
  OA22X1 U4645 ( .IN1(n6271), .IN2(n5361), .IN3(n5353), .IN4(n6117), .Q(n3863)
         );
  OAI22X1 U4646 ( .IN1(n6426), .IN2(n5404), .IN3(n5403), .IN4(n3864), .QN(
        N10254) );
  OA22X1 U4647 ( .IN1(n6426), .IN2(n5381), .IN3(n5389), .IN4(n3865), .Q(n3864)
         );
  OA22X1 U4648 ( .IN1(n5371), .IN2(n3866), .IN3(n6272), .IN4(n5366), .Q(n3865)
         );
  OA22X1 U4649 ( .IN1(n6272), .IN2(n5361), .IN3(n5353), .IN4(n6118), .Q(n3866)
         );
  OAI22X1 U4650 ( .IN1(n6427), .IN2(n5397), .IN3(n5403), .IN4(n3867), .QN(
        N10253) );
  OA22X1 U4651 ( .IN1(n6427), .IN2(n5381), .IN3(n5395), .IN4(n3868), .Q(n3867)
         );
  OA22X1 U4652 ( .IN1(n5371), .IN2(n3869), .IN3(n6273), .IN4(n5366), .Q(n3868)
         );
  OA22X1 U4653 ( .IN1(n6273), .IN2(n5362), .IN3(n5353), .IN4(n6119), .Q(n3869)
         );
  OAI22X1 U4654 ( .IN1(n6428), .IN2(n5406), .IN3(n5403), .IN4(n3870), .QN(
        N10252) );
  OA22X1 U4655 ( .IN1(n6428), .IN2(n5381), .IN3(n5394), .IN4(n3871), .Q(n3870)
         );
  OA22X1 U4656 ( .IN1(n5371), .IN2(n3872), .IN3(n6274), .IN4(n5366), .Q(n3871)
         );
  OA22X1 U4657 ( .IN1(n6274), .IN2(n5362), .IN3(n5353), .IN4(n6120), .Q(n3872)
         );
  OAI22X1 U4658 ( .IN1(n6429), .IN2(n5405), .IN3(n5403), .IN4(n3873), .QN(
        N10251) );
  OA22X1 U4659 ( .IN1(n6429), .IN2(n5381), .IN3(n5396), .IN4(n3874), .Q(n3873)
         );
  OA22X1 U4660 ( .IN1(n5371), .IN2(n3875), .IN3(n6275), .IN4(n5366), .Q(n3874)
         );
  OA22X1 U4661 ( .IN1(n6275), .IN2(n5362), .IN3(n5353), .IN4(n6121), .Q(n3875)
         );
  OAI22X1 U4662 ( .IN1(n6430), .IN2(n5397), .IN3(n5403), .IN4(n3876), .QN(
        N10250) );
  OA22X1 U4663 ( .IN1(n6430), .IN2(n5381), .IN3(n5391), .IN4(n3877), .Q(n3876)
         );
  OA22X1 U4664 ( .IN1(n5371), .IN2(n3878), .IN3(n6276), .IN4(n5366), .Q(n3877)
         );
  OA22X1 U4665 ( .IN1(n6276), .IN2(n5362), .IN3(n5353), .IN4(n6122), .Q(n3878)
         );
  OAI22X1 U4666 ( .IN1(n6431), .IN2(n5404), .IN3(n5403), .IN4(n3879), .QN(
        N10249) );
  OA22X1 U4667 ( .IN1(n6431), .IN2(n5381), .IN3(n5391), .IN4(n3880), .Q(n3879)
         );
  OA22X1 U4668 ( .IN1(n5371), .IN2(n3881), .IN3(n6277), .IN4(n5366), .Q(n3880)
         );
  OA22X1 U4669 ( .IN1(n6277), .IN2(n5362), .IN3(n5353), .IN4(n6123), .Q(n3881)
         );
  OAI22X1 U4670 ( .IN1(n6432), .IN2(n5405), .IN3(n5403), .IN4(n3882), .QN(
        N10248) );
  OA22X1 U4671 ( .IN1(n6432), .IN2(n5381), .IN3(n5388), .IN4(n3883), .Q(n3882)
         );
  OA22X1 U4672 ( .IN1(n5371), .IN2(n3884), .IN3(n6278), .IN4(n5366), .Q(n3883)
         );
  OA22X1 U4673 ( .IN1(n6278), .IN2(n5361), .IN3(n5353), .IN4(n6124), .Q(n3884)
         );
  OAI22X1 U4674 ( .IN1(n6433), .IN2(n5406), .IN3(n5403), .IN4(n3885), .QN(
        N10247) );
  OA22X1 U4675 ( .IN1(n6433), .IN2(n5381), .IN3(n5390), .IN4(n3886), .Q(n3885)
         );
  OA22X1 U4676 ( .IN1(n5371), .IN2(n3887), .IN3(n6279), .IN4(n5366), .Q(n3886)
         );
  OA22X1 U4677 ( .IN1(n6279), .IN2(n5356), .IN3(n5353), .IN4(n6125), .Q(n3887)
         );
  OAI22X1 U4678 ( .IN1(n6434), .IN2(n5408), .IN3(n5403), .IN4(n3888), .QN(
        N10246) );
  OA22X1 U4679 ( .IN1(n6434), .IN2(n5381), .IN3(n5386), .IN4(n3889), .Q(n3888)
         );
  OA22X1 U4680 ( .IN1(n5371), .IN2(n3890), .IN3(n6280), .IN4(n5366), .Q(n3889)
         );
  OA22X1 U4681 ( .IN1(n6280), .IN2(n5357), .IN3(n5353), .IN4(n6126), .Q(n3890)
         );
  OAI22X1 U4682 ( .IN1(n6435), .IN2(n5398), .IN3(n5403), .IN4(n3891), .QN(
        N10245) );
  OA22X1 U4683 ( .IN1(n6435), .IN2(n5381), .IN3(n5387), .IN4(n3892), .Q(n3891)
         );
  OA22X1 U4684 ( .IN1(n5371), .IN2(n3893), .IN3(n6281), .IN4(n5366), .Q(n3892)
         );
  OA22X1 U4685 ( .IN1(n6281), .IN2(n5358), .IN3(n5353), .IN4(n6127), .Q(n3893)
         );
  OAI22X1 U4686 ( .IN1(n6436), .IN2(n5397), .IN3(n5403), .IN4(n3894), .QN(
        N10244) );
  OA22X1 U4687 ( .IN1(n6436), .IN2(n5381), .IN3(n5386), .IN4(n3895), .Q(n3894)
         );
  OA22X1 U4688 ( .IN1(n5370), .IN2(n3896), .IN3(n6282), .IN4(n5366), .Q(n3895)
         );
  OA22X1 U4689 ( .IN1(n6282), .IN2(n5357), .IN3(n5353), .IN4(n6128), .Q(n3896)
         );
  OAI22X1 U4690 ( .IN1(n6437), .IN2(n5409), .IN3(n5403), .IN4(n3897), .QN(
        N10243) );
  OA22X1 U4691 ( .IN1(n6437), .IN2(n5380), .IN3(n5386), .IN4(n3898), .Q(n3897)
         );
  OA22X1 U4692 ( .IN1(n5370), .IN2(n3899), .IN3(n6283), .IN4(n5366), .Q(n3898)
         );
  OA22X1 U4693 ( .IN1(n6283), .IN2(n5357), .IN3(n5353), .IN4(n6129), .Q(n3899)
         );
  OAI22X1 U4694 ( .IN1(n6438), .IN2(n5407), .IN3(n5403), .IN4(n3900), .QN(
        N10242) );
  OA22X1 U4695 ( .IN1(n6438), .IN2(n5380), .IN3(n5386), .IN4(n3901), .Q(n3900)
         );
  OA22X1 U4696 ( .IN1(n5370), .IN2(n3902), .IN3(n6284), .IN4(n5366), .Q(n3901)
         );
  OA22X1 U4697 ( .IN1(n6284), .IN2(n5358), .IN3(n5353), .IN4(n6130), .Q(n3902)
         );
  OAI22X1 U4698 ( .IN1(n6439), .IN2(n5406), .IN3(n5403), .IN4(n3903), .QN(
        N10241) );
  OA22X1 U4699 ( .IN1(n6439), .IN2(n5380), .IN3(n5386), .IN4(n3904), .Q(n3903)
         );
  OA22X1 U4700 ( .IN1(n5370), .IN2(n3905), .IN3(n6285), .IN4(n5366), .Q(n3904)
         );
  OA22X1 U4701 ( .IN1(n6285), .IN2(n5359), .IN3(n5353), .IN4(n6131), .Q(n3905)
         );
  OAI22X1 U4702 ( .IN1(n6440), .IN2(n5397), .IN3(n5403), .IN4(n3906), .QN(
        N10240) );
  OA22X1 U4703 ( .IN1(n6440), .IN2(n5380), .IN3(n5386), .IN4(n3907), .Q(n3906)
         );
  OA22X1 U4704 ( .IN1(n5370), .IN2(n3908), .IN3(n6286), .IN4(n5366), .Q(n3907)
         );
  OA22X1 U4705 ( .IN1(n6286), .IN2(n5360), .IN3(n5353), .IN4(n6132), .Q(n3908)
         );
  OAI22X1 U4706 ( .IN1(n6441), .IN2(n5408), .IN3(n5403), .IN4(n3909), .QN(
        N10239) );
  OA22X1 U4707 ( .IN1(n6441), .IN2(n5380), .IN3(n5387), .IN4(n3910), .Q(n3909)
         );
  OA22X1 U4708 ( .IN1(n5370), .IN2(n3911), .IN3(n6287), .IN4(n5366), .Q(n3910)
         );
  OA22X1 U4709 ( .IN1(n6287), .IN2(n5358), .IN3(n5353), .IN4(n6133), .Q(n3911)
         );
  OAI22X1 U4710 ( .IN1(n6442), .IN2(n5397), .IN3(n5403), .IN4(n3912), .QN(
        N10238) );
  OA22X1 U4711 ( .IN1(n6442), .IN2(n5380), .IN3(n5387), .IN4(n3913), .Q(n3912)
         );
  OA22X1 U4712 ( .IN1(n5370), .IN2(n3914), .IN3(n6288), .IN4(n5366), .Q(n3913)
         );
  OA22X1 U4713 ( .IN1(n6288), .IN2(n5362), .IN3(n5269), .IN4(n6134), .Q(n3914)
         );
  OAI22X1 U4714 ( .IN1(n6443), .IN2(n5409), .IN3(n5403), .IN4(n3915), .QN(
        N10236) );
  OA22X1 U4715 ( .IN1(n6443), .IN2(n5380), .IN3(n5387), .IN4(n3916), .Q(n3915)
         );
  OA22X1 U4716 ( .IN1(n5370), .IN2(n3917), .IN3(n6289), .IN4(n5366), .Q(n3916)
         );
  OA22X1 U4717 ( .IN1(n6289), .IN2(n5359), .IN3(n5269), .IN4(n6135), .Q(n3917)
         );
  OAI22X1 U4718 ( .IN1(n6444), .IN2(n5398), .IN3(n5403), .IN4(n3918), .QN(
        N10235) );
  OA22X1 U4719 ( .IN1(n6444), .IN2(n5380), .IN3(n5387), .IN4(n3919), .Q(n3918)
         );
  OA22X1 U4720 ( .IN1(n5370), .IN2(n3920), .IN3(n6290), .IN4(n5366), .Q(n3919)
         );
  OA22X1 U4721 ( .IN1(n6290), .IN2(n5361), .IN3(n5269), .IN4(n6136), .Q(n3920)
         );
  OAI22X1 U4722 ( .IN1(n6445), .IN2(n5404), .IN3(n5403), .IN4(n3921), .QN(
        N10234) );
  OA22X1 U4723 ( .IN1(n6445), .IN2(n5380), .IN3(n5387), .IN4(n3922), .Q(n3921)
         );
  OA22X1 U4724 ( .IN1(n5370), .IN2(n3923), .IN3(n6291), .IN4(n5366), .Q(n3922)
         );
  OA22X1 U4725 ( .IN1(n6291), .IN2(n5355), .IN3(n5269), .IN4(n6137), .Q(n3923)
         );
  OAI22X1 U4726 ( .IN1(n6446), .IN2(n5405), .IN3(n5403), .IN4(n3924), .QN(
        N10233) );
  OA22X1 U4727 ( .IN1(n6446), .IN2(n5380), .IN3(n5388), .IN4(n3925), .Q(n3924)
         );
  OA22X1 U4728 ( .IN1(n5370), .IN2(n3926), .IN3(n6292), .IN4(n5366), .Q(n3925)
         );
  OA22X1 U4729 ( .IN1(n6292), .IN2(n5358), .IN3(n5269), .IN4(n6138), .Q(n3926)
         );
  OAI22X1 U4730 ( .IN1(n6447), .IN2(n5406), .IN3(n5403), .IN4(n3927), .QN(
        N10232) );
  OA22X1 U4731 ( .IN1(n6447), .IN2(n5380), .IN3(n5388), .IN4(n3928), .Q(n3927)
         );
  OA22X1 U4732 ( .IN1(n5370), .IN2(n3929), .IN3(n6293), .IN4(n5366), .Q(n3928)
         );
  OA22X1 U4733 ( .IN1(n6293), .IN2(n5359), .IN3(n5269), .IN4(n6139), .Q(n3929)
         );
  OAI22X1 U4734 ( .IN1(n6448), .IN2(n5398), .IN3(n5403), .IN4(n3930), .QN(
        N10231) );
  OA22X1 U4735 ( .IN1(n6448), .IN2(n5380), .IN3(n5388), .IN4(n3931), .Q(n3930)
         );
  OA22X1 U4736 ( .IN1(n5369), .IN2(n3932), .IN3(n6294), .IN4(n5366), .Q(n3931)
         );
  OA22X1 U4737 ( .IN1(n6294), .IN2(n5360), .IN3(n5269), .IN4(n6140), .Q(n3932)
         );
  OAI22X1 U4738 ( .IN1(n6449), .IN2(n5398), .IN3(n5403), .IN4(n3933), .QN(
        N10230) );
  OA22X1 U4739 ( .IN1(n6449), .IN2(n5380), .IN3(n5388), .IN4(n3934), .Q(n3933)
         );
  OA22X1 U4740 ( .IN1(n5369), .IN2(n3935), .IN3(n6295), .IN4(n5366), .Q(n3934)
         );
  OA22X1 U4741 ( .IN1(n6295), .IN2(n5361), .IN3(n5269), .IN4(n6141), .Q(n3935)
         );
  OAI22X1 U4742 ( .IN1(n6450), .IN2(n5397), .IN3(n5403), .IN4(n3936), .QN(
        N10229) );
  OA22X1 U4743 ( .IN1(n6450), .IN2(n5380), .IN3(n5388), .IN4(n3937), .Q(n3936)
         );
  OA22X1 U4744 ( .IN1(n5369), .IN2(n3938), .IN3(n6296), .IN4(n5366), .Q(n3937)
         );
  OA22X1 U4745 ( .IN1(n6296), .IN2(n5359), .IN3(n5269), .IN4(n6142), .Q(n3938)
         );
  OAI22X1 U4746 ( .IN1(n6451), .IN2(n5405), .IN3(n5403), .IN4(n3939), .QN(
        N10228) );
  OA22X1 U4747 ( .IN1(n6451), .IN2(n5379), .IN3(n5389), .IN4(n3940), .Q(n3939)
         );
  OA22X1 U4748 ( .IN1(n5369), .IN2(n3941), .IN3(n6297), .IN4(n5366), .Q(n3940)
         );
  OA22X1 U4749 ( .IN1(n6297), .IN2(n5361), .IN3(n5269), .IN4(n6143), .Q(n3941)
         );
  OAI22X1 U4750 ( .IN1(n6452), .IN2(n5408), .IN3(n5403), .IN4(n3942), .QN(
        N10227) );
  OA22X1 U4751 ( .IN1(n6452), .IN2(n5379), .IN3(n5389), .IN4(n3943), .Q(n3942)
         );
  OA22X1 U4752 ( .IN1(n5369), .IN2(n3944), .IN3(n6298), .IN4(n5366), .Q(n3943)
         );
  OA22X1 U4753 ( .IN1(n6298), .IN2(n5355), .IN3(n5269), .IN4(n6144), .Q(n3944)
         );
  OAI22X1 U4754 ( .IN1(n6453), .IN2(n5398), .IN3(n5403), .IN4(n3945), .QN(
        N10226) );
  OA22X1 U4755 ( .IN1(n6453), .IN2(n5379), .IN3(n5389), .IN4(n3946), .Q(n3945)
         );
  OA22X1 U4756 ( .IN1(n5369), .IN2(n3947), .IN3(n6299), .IN4(n5366), .Q(n3946)
         );
  OA22X1 U4757 ( .IN1(n6299), .IN2(n5356), .IN3(n5269), .IN4(n6145), .Q(n3947)
         );
  OAI22X1 U4758 ( .IN1(n6454), .IN2(n5406), .IN3(n5400), .IN4(n3948), .QN(
        N10225) );
  OA22X1 U4759 ( .IN1(n6454), .IN2(n5379), .IN3(n5389), .IN4(n3949), .Q(n3948)
         );
  OA22X1 U4760 ( .IN1(n5369), .IN2(n3950), .IN3(n6300), .IN4(n5366), .Q(n3949)
         );
  OA22X1 U4761 ( .IN1(n6300), .IN2(n5357), .IN3(n5269), .IN4(n6146), .Q(n3950)
         );
  OA22X1 U4763 ( .IN1(n6320), .IN2(n5379), .IN3(n5389), .IN4(n3952), .Q(n3951)
         );
  OA22X1 U4767 ( .IN1(n6321), .IN2(n5379), .IN3(n5390), .IN4(n3955), .Q(n3954)
         );
  OA22X1 U4771 ( .IN1(n6322), .IN2(n5379), .IN3(n5390), .IN4(n3958), .Q(n3957)
         );
  OA22X1 U4775 ( .IN1(n6323), .IN2(n5379), .IN3(n5390), .IN4(n3961), .Q(n3960)
         );
  OA22X1 U4779 ( .IN1(n6324), .IN2(n5379), .IN3(n5390), .IN4(n3964), .Q(n3963)
         );
  OA22X1 U4783 ( .IN1(n6325), .IN2(n5379), .IN3(n5390), .IN4(n3967), .Q(n3966)
         );
  OA22X1 U4787 ( .IN1(n6326), .IN2(n5379), .IN3(n5391), .IN4(n3970), .Q(n3969)
         );
  OA22X1 U4791 ( .IN1(n6327), .IN2(n5379), .IN3(n5391), .IN4(n3973), .Q(n3972)
         );
  OA22X1 U4795 ( .IN1(n6328), .IN2(n5379), .IN3(n5391), .IN4(n3976), .Q(n3975)
         );
  OA22X1 U4799 ( .IN1(n6329), .IN2(n5379), .IN3(n5391), .IN4(n3979), .Q(n3978)
         );
  OA22X1 U4803 ( .IN1(n6330), .IN2(n5378), .IN3(n5391), .IN4(n3982), .Q(n3981)
         );
  OA22X1 U4807 ( .IN1(n6331), .IN2(n5378), .IN3(n5392), .IN4(n3985), .Q(n3984)
         );
  OA22X1 U4811 ( .IN1(n6332), .IN2(n5378), .IN3(n5392), .IN4(n3988), .Q(n3987)
         );
  OA22X1 U4815 ( .IN1(n6333), .IN2(n5378), .IN3(n5392), .IN4(n3991), .Q(n3990)
         );
  OA22X1 U4819 ( .IN1(n6334), .IN2(n5378), .IN3(n5392), .IN4(n3994), .Q(n3993)
         );
  OA22X1 U4823 ( .IN1(n6335), .IN2(n5378), .IN3(n5392), .IN4(n3997), .Q(n3996)
         );
  OA22X1 U4827 ( .IN1(n6336), .IN2(n5378), .IN3(n5393), .IN4(n4000), .Q(n3999)
         );
  OA22X1 U4831 ( .IN1(n6337), .IN2(n5378), .IN3(n5393), .IN4(n4003), .Q(n4002)
         );
  OA22X1 U4835 ( .IN1(n6338), .IN2(n5378), .IN3(n5393), .IN4(n4006), .Q(n4005)
         );
  OA22X1 U4839 ( .IN1(n6339), .IN2(n5378), .IN3(n5393), .IN4(n4009), .Q(n4008)
         );
  OA22X1 U4843 ( .IN1(n6340), .IN2(n5378), .IN3(n5393), .IN4(n4012), .Q(n4011)
         );
  OA22X1 U4847 ( .IN1(n6341), .IN2(n5378), .IN3(n5389), .IN4(n4015), .Q(n4014)
         );
  OA22X1 U4851 ( .IN1(n6342), .IN2(n5378), .IN3(n5394), .IN4(n4018), .Q(n4017)
         );
  OA22X1 U4855 ( .IN1(n6343), .IN2(n5378), .IN3(n5395), .IN4(n4021), .Q(n4020)
         );
  OA22X1 U4859 ( .IN1(n6344), .IN2(n5377), .IN3(n5391), .IN4(n4024), .Q(n4023)
         );
  OA22X1 U4863 ( .IN1(n6345), .IN2(n5377), .IN3(n5388), .IN4(n4027), .Q(n4026)
         );
  OA22X1 U4867 ( .IN1(n6346), .IN2(n5377), .IN3(n5390), .IN4(n4030), .Q(n4029)
         );
  OA22X1 U4871 ( .IN1(n6315), .IN2(n5377), .IN3(n5391), .IN4(n4033), .Q(n4032)
         );
  OA22X1 U4875 ( .IN1(n6316), .IN2(n5377), .IN3(n5386), .IN4(n4036), .Q(n4035)
         );
  OA22X1 U4879 ( .IN1(n6317), .IN2(n5377), .IN3(n5387), .IN4(n4039), .Q(n4038)
         );
  OA22X1 U4883 ( .IN1(n6318), .IN2(n5377), .IN3(n5388), .IN4(n4042), .Q(n4041)
         );
  OA22X1 U4887 ( .IN1(n6319), .IN2(n5377), .IN3(n5393), .IN4(n4045), .Q(n4044)
         );
  OAI22X1 U4890 ( .IN1(n6455), .IN2(n5397), .IN3(n5399), .IN4(n4047), .QN(
        N10192) );
  OA22X1 U4891 ( .IN1(n6455), .IN2(n5377), .IN3(n5392), .IN4(n4048), .Q(n4047)
         );
  OA22X1 U4892 ( .IN1(n5369), .IN2(n4049), .IN3(n6301), .IN4(n5365), .Q(n4048)
         );
  OA22X1 U4893 ( .IN1(n6301), .IN2(n5362), .IN3(n5269), .IN4(n6147), .Q(n4049)
         );
  OAI22X1 U4894 ( .IN1(n6456), .IN2(n5397), .IN3(n5400), .IN4(n4050), .QN(
        N10191) );
  OA22X1 U4895 ( .IN1(n6456), .IN2(n5377), .IN3(n5390), .IN4(n4051), .Q(n4050)
         );
  OA22X1 U4896 ( .IN1(n5369), .IN2(n4052), .IN3(n6302), .IN4(n5365), .Q(n4051)
         );
  OA22X1 U4897 ( .IN1(n6302), .IN2(n5362), .IN3(n5269), .IN4(n6148), .Q(n4052)
         );
  OAI22X1 U4898 ( .IN1(n6457), .IN2(n5397), .IN3(n5399), .IN4(n4053), .QN(
        N10190) );
  OA22X1 U4899 ( .IN1(n6457), .IN2(n5377), .IN3(n5390), .IN4(n4054), .Q(n4053)
         );
  OA22X1 U4900 ( .IN1(n5369), .IN2(n4055), .IN3(n6303), .IN4(n5365), .Q(n4054)
         );
  OA22X1 U4901 ( .IN1(n6303), .IN2(n5362), .IN3(n5269), .IN4(n6149), .Q(n4055)
         );
  OAI22X1 U4902 ( .IN1(n6458), .IN2(n5408), .IN3(n5400), .IN4(n4056), .QN(
        N10189) );
  OA22X1 U4903 ( .IN1(n6458), .IN2(n5377), .IN3(n5394), .IN4(n4057), .Q(n4056)
         );
  OA22X1 U4904 ( .IN1(n5369), .IN2(n4058), .IN3(n6304), .IN4(n5365), .Q(n4057)
         );
  OA22X1 U4905 ( .IN1(n6304), .IN2(n5358), .IN3(n5269), .IN4(n6150), .Q(n4058)
         );
  OAI22X1 U4906 ( .IN1(n6459), .IN2(n5405), .IN3(n5399), .IN4(n4059), .QN(
        N10188) );
  OA22X1 U4907 ( .IN1(n6459), .IN2(n5377), .IN3(n5394), .IN4(n4060), .Q(n4059)
         );
  OA22X1 U4908 ( .IN1(n5369), .IN2(n4061), .IN3(n6305), .IN4(n5365), .Q(n4060)
         );
  OA22X1 U4909 ( .IN1(n6305), .IN2(n5359), .IN3(n5353), .IN4(n6151), .Q(n4061)
         );
  NAND4X0 U4910 ( .IN1(n4062), .IN2(n5377), .IN3(n4063), .IN4(n5365), .QN(
        decodedVector_o[4]) );
  NAND4X0 U4912 ( .IN1(decodedPacketValid[4]), .IN2(n2908), .IN3(n5995), .IN4(
        n5990), .QN(n3686) );
  NAND4X0 U4913 ( .IN1(decodedPacketValid[7]), .IN2(n2909), .IN3(n5992), .IN4(
        n5987), .QN(n3680) );
  NAND4X0 U4914 ( .IN1(decodedPacketValid[6]), .IN2(n2910), .IN3(n5993), .IN4(
        n5988), .QN(n3682) );
  NAND4X0 U4915 ( .IN1(decodedPacketValid[3]), .IN2(N1070), .IN3(n5996), .IN4(
        n5991), .QN(n4062) );
  OA22X1 U4937 ( .IN1(n5321), .IN2(n4091), .IN3(n5856), .IN4(n5334), .Q(n4090)
         );
  OAI22X1 U4941 ( .IN1(n5340), .IN2(n4094), .IN3(n6384), .IN4(n5343), .QN(
        N10181) );
  OA22X1 U4942 ( .IN1(n5321), .IN2(n4095), .IN3(n6349), .IN4(n5319), .Q(n4094)
         );
  OA22X1 U4943 ( .IN1(n6230), .IN2(n5309), .IN3(n5317), .IN4(n4096), .Q(n4095)
         );
  OA22X1 U4944 ( .IN1(n5286), .IN2(n4097), .IN3(n6195), .IN4(n5296), .Q(n4096)
         );
  OA22X1 U4945 ( .IN1(n6076), .IN2(n5281), .IN3(n5282), .IN4(n6041), .Q(n4097)
         );
  OAI22X1 U4946 ( .IN1(n5340), .IN2(n4098), .IN3(n6376), .IN4(n5349), .QN(
        N10180) );
  OA22X1 U4947 ( .IN1(n5321), .IN2(n4099), .IN3(n6348), .IN4(n5331), .Q(n4098)
         );
  OA22X1 U4948 ( .IN1(n6222), .IN2(n5309), .IN3(n5314), .IN4(n4100), .Q(n4099)
         );
  OA22X1 U4949 ( .IN1(n5286), .IN2(n4101), .IN3(n6194), .IN4(n5296), .Q(n4100)
         );
  OA22X1 U4950 ( .IN1(n6068), .IN2(n5281), .IN3(n5283), .IN4(n6040), .Q(n4101)
         );
  OAI22X1 U4951 ( .IN1(n5340), .IN2(n4102), .IN3(n6372), .IN4(n5344), .QN(
        N10179) );
  OA22X1 U4952 ( .IN1(n5321), .IN2(n4103), .IN3(n6374), .IN4(n5331), .Q(n4102)
         );
  OA22X1 U4953 ( .IN1(n6218), .IN2(n5309), .IN3(n5317), .IN4(n4104), .Q(n4103)
         );
  OA22X1 U4954 ( .IN1(n5286), .IN2(n4105), .IN3(n6220), .IN4(n5297), .Q(n4104)
         );
  OA22X1 U4955 ( .IN1(n6064), .IN2(n5281), .IN3(n5283), .IN4(n6066), .Q(n4105)
         );
  OA22X1 U4957 ( .IN1(n5321), .IN2(n4107), .IN3(n6371), .IN4(n5331), .Q(n4106)
         );
  OAI22X1 U4961 ( .IN1(n5340), .IN2(n4110), .IN3(n6373), .IN4(n5345), .QN(
        N10177) );
  OA22X1 U4962 ( .IN1(n5321), .IN2(n4111), .IN3(n6370), .IN4(n5331), .Q(n4110)
         );
  OA22X1 U4963 ( .IN1(n6219), .IN2(n5309), .IN3(n5313), .IN4(n4112), .Q(n4111)
         );
  OA22X1 U4964 ( .IN1(n5286), .IN2(n4113), .IN3(n6216), .IN4(n5297), .Q(n4112)
         );
  OA22X1 U4965 ( .IN1(n6065), .IN2(n5281), .IN3(n5283), .IN4(n6062), .Q(n4113)
         );
  OAI22X1 U4966 ( .IN1(n5341), .IN2(n4114), .IN3(n6398), .IN4(n5346), .QN(
        N10176) );
  OA22X1 U4967 ( .IN1(n5321), .IN2(n4115), .IN3(n6347), .IN4(n5331), .Q(n4114)
         );
  OA22X1 U4968 ( .IN1(n6245), .IN2(n5309), .IN3(n5310), .IN4(n4116), .Q(n4115)
         );
  OA22X1 U4969 ( .IN1(n5286), .IN2(n4117), .IN3(n6193), .IN4(n5297), .Q(n4116)
         );
  OA22X1 U4970 ( .IN1(n6091), .IN2(n5281), .IN3(n5283), .IN4(n6039), .Q(n4117)
         );
  OAI22X1 U4971 ( .IN1(n5341), .IN2(n4118), .IN3(n5967), .IN4(n5350), .QN(
        N10175) );
  OA22X1 U4972 ( .IN1(n5321), .IN2(n4119), .IN3(n6369), .IN4(n5331), .Q(n4118)
         );
  OA22X1 U4973 ( .IN1(n5952), .IN2(n5309), .IN3(n5310), .IN4(n4120), .Q(n4119)
         );
  OA22X1 U4974 ( .IN1(n5286), .IN2(n4121), .IN3(n6215), .IN4(n5297), .Q(n4120)
         );
  OA22X1 U4975 ( .IN1(n5937), .IN2(n5281), .IN3(n5283), .IN4(n6061), .Q(n4121)
         );
  OAI22X1 U4976 ( .IN1(n5341), .IN2(n4122), .IN3(n5968), .IN4(n5345), .QN(
        N10174) );
  OA22X1 U4977 ( .IN1(n5321), .IN2(n4123), .IN3(n6368), .IN4(n5331), .Q(n4122)
         );
  OA22X1 U4978 ( .IN1(n5953), .IN2(n5309), .IN3(n5310), .IN4(n4124), .Q(n4123)
         );
  OA22X1 U4979 ( .IN1(n5286), .IN2(n4125), .IN3(n6214), .IN4(n5297), .Q(n4124)
         );
  OA22X1 U4980 ( .IN1(n5938), .IN2(n5281), .IN3(n5283), .IN4(n6060), .Q(n4125)
         );
  OAI22X1 U4981 ( .IN1(n5341), .IN2(n4126), .IN3(n5969), .IN4(n5348), .QN(
        N10173) );
  OA22X1 U4982 ( .IN1(n5321), .IN2(n4127), .IN3(n6367), .IN4(n5331), .Q(n4126)
         );
  OA22X1 U4983 ( .IN1(n5954), .IN2(n5309), .IN3(n5310), .IN4(n4128), .Q(n4127)
         );
  OA22X1 U4984 ( .IN1(n5286), .IN2(n4129), .IN3(n6213), .IN4(n5297), .Q(n4128)
         );
  OA22X1 U4985 ( .IN1(n5939), .IN2(n5281), .IN3(n5283), .IN4(n6059), .Q(n4129)
         );
  OAI22X1 U4986 ( .IN1(n5341), .IN2(n4130), .IN3(n5970), .IN4(n5350), .QN(
        N10172) );
  OA22X1 U4987 ( .IN1(n5321), .IN2(n4131), .IN3(n6366), .IN4(n5331), .Q(n4130)
         );
  OA22X1 U4988 ( .IN1(n5955), .IN2(n5309), .IN3(n5310), .IN4(n4132), .Q(n4131)
         );
  OA22X1 U4989 ( .IN1(n5286), .IN2(n4133), .IN3(n6212), .IN4(n5297), .Q(n4132)
         );
  OA22X1 U4990 ( .IN1(n5940), .IN2(n5281), .IN3(n5283), .IN4(n6058), .Q(n4133)
         );
  OAI22X1 U4991 ( .IN1(n5341), .IN2(n4134), .IN3(n5971), .IN4(n5349), .QN(
        N10171) );
  OA22X1 U4992 ( .IN1(n5321), .IN2(n4135), .IN3(n6365), .IN4(n5331), .Q(n4134)
         );
  OA22X1 U4993 ( .IN1(n5956), .IN2(n5309), .IN3(n5311), .IN4(n4136), .Q(n4135)
         );
  OA22X1 U4994 ( .IN1(n5286), .IN2(n4137), .IN3(n6211), .IN4(n5297), .Q(n4136)
         );
  OA22X1 U4995 ( .IN1(n5941), .IN2(n5281), .IN3(n5283), .IN4(n6057), .Q(n4137)
         );
  OAI22X1 U4996 ( .IN1(n5341), .IN2(n4138), .IN3(n5972), .IN4(n5347), .QN(
        N10170) );
  OA22X1 U4997 ( .IN1(n5322), .IN2(n4139), .IN3(n6364), .IN4(n5331), .Q(n4138)
         );
  OA22X1 U4998 ( .IN1(n5957), .IN2(n5309), .IN3(n5314), .IN4(n4140), .Q(n4139)
         );
  OA22X1 U4999 ( .IN1(n5287), .IN2(n4141), .IN3(n6210), .IN4(n5297), .Q(n4140)
         );
  OA22X1 U5000 ( .IN1(n5942), .IN2(n5281), .IN3(n5283), .IN4(n6056), .Q(n4141)
         );
  OAI22X1 U5001 ( .IN1(n5341), .IN2(n4142), .IN3(n5973), .IN4(n5349), .QN(
        N10169) );
  OA22X1 U5002 ( .IN1(n5322), .IN2(n4143), .IN3(n6363), .IN4(n5331), .Q(n4142)
         );
  OA22X1 U5003 ( .IN1(n5958), .IN2(n5309), .IN3(n5314), .IN4(n4144), .Q(n4143)
         );
  OA22X1 U5004 ( .IN1(n5287), .IN2(n4145), .IN3(n6209), .IN4(n5297), .Q(n4144)
         );
  OA22X1 U5005 ( .IN1(n5943), .IN2(n5281), .IN3(n5283), .IN4(n6055), .Q(n4145)
         );
  OAI22X1 U5006 ( .IN1(n5341), .IN2(n4146), .IN3(n5974), .IN4(n5348), .QN(
        N10168) );
  OA22X1 U5007 ( .IN1(n5322), .IN2(n4147), .IN3(n6362), .IN4(n5331), .Q(n4146)
         );
  OA22X1 U5008 ( .IN1(n5959), .IN2(n5309), .IN3(n5314), .IN4(n4148), .Q(n4147)
         );
  OA22X1 U5009 ( .IN1(n5287), .IN2(n4149), .IN3(n6208), .IN4(n5297), .Q(n4148)
         );
  OA22X1 U5010 ( .IN1(n5944), .IN2(n5281), .IN3(n5283), .IN4(n6054), .Q(n4149)
         );
  OAI22X1 U5011 ( .IN1(n5341), .IN2(n4150), .IN3(n5975), .IN4(n5349), .QN(
        N10167) );
  OA22X1 U5012 ( .IN1(n5322), .IN2(n4151), .IN3(n6308), .IN4(n5331), .Q(n4150)
         );
  OA22X1 U5013 ( .IN1(n5960), .IN2(n5309), .IN3(n5317), .IN4(n4152), .Q(n4151)
         );
  OA22X1 U5014 ( .IN1(n5287), .IN2(n4153), .IN3(n6154), .IN4(n5297), .Q(n4152)
         );
  OA22X1 U5015 ( .IN1(n5945), .IN2(n5281), .IN3(n5283), .IN4(n6000), .Q(n4153)
         );
  OAI22X1 U5016 ( .IN1(n5341), .IN2(n4154), .IN3(n5976), .IN4(n5343), .QN(
        N10166) );
  OA22X1 U5017 ( .IN1(n5322), .IN2(n4155), .IN3(n6309), .IN4(n5331), .Q(n4154)
         );
  OA22X1 U5018 ( .IN1(n5961), .IN2(n5309), .IN3(n5312), .IN4(n4156), .Q(n4155)
         );
  OA22X1 U5019 ( .IN1(n5287), .IN2(n4157), .IN3(n6155), .IN4(n5297), .Q(n4156)
         );
  OA22X1 U5020 ( .IN1(n5946), .IN2(n5281), .IN3(n5283), .IN4(n6001), .Q(n4157)
         );
  OAI22X1 U5021 ( .IN1(n5341), .IN2(n4158), .IN3(n5977), .IN4(n5343), .QN(
        N10165) );
  OA22X1 U5022 ( .IN1(n5322), .IN2(n4159), .IN3(n6310), .IN4(n5332), .Q(n4158)
         );
  OA22X1 U5023 ( .IN1(n5962), .IN2(n5309), .IN3(n5314), .IN4(n4160), .Q(n4159)
         );
  OA22X1 U5024 ( .IN1(n5287), .IN2(n4161), .IN3(n6156), .IN4(n5297), .Q(n4160)
         );
  OA22X1 U5025 ( .IN1(n5947), .IN2(n5281), .IN3(n5283), .IN4(n6002), .Q(n4161)
         );
  OAI22X1 U5026 ( .IN1(n5341), .IN2(n4162), .IN3(n5978), .IN4(n5350), .QN(
        N10164) );
  OA22X1 U5027 ( .IN1(n5322), .IN2(n4163), .IN3(n6311), .IN4(n5332), .Q(n4162)
         );
  OA22X1 U5028 ( .IN1(n5963), .IN2(n5309), .IN3(n5317), .IN4(n4164), .Q(n4163)
         );
  OA22X1 U5029 ( .IN1(n5287), .IN2(n4165), .IN3(n6157), .IN4(n5298), .Q(n4164)
         );
  OA22X1 U5030 ( .IN1(n5948), .IN2(n5280), .IN3(n5283), .IN4(n6003), .Q(n4165)
         );
  OAI22X1 U5031 ( .IN1(n5341), .IN2(n4166), .IN3(n5979), .IN4(n5350), .QN(
        N10163) );
  OA22X1 U5032 ( .IN1(n5322), .IN2(n4167), .IN3(n6312), .IN4(n5332), .Q(n4166)
         );
  OA22X1 U5033 ( .IN1(n5964), .IN2(n5308), .IN3(n5312), .IN4(n4168), .Q(n4167)
         );
  OA22X1 U5034 ( .IN1(n5287), .IN2(n4169), .IN3(n6158), .IN4(n5298), .Q(n4168)
         );
  OA22X1 U5035 ( .IN1(n5949), .IN2(n5280), .IN3(n5283), .IN4(n6004), .Q(n4169)
         );
  OAI22X1 U5036 ( .IN1(n5341), .IN2(n4170), .IN3(n5980), .IN4(n5349), .QN(
        N10162) );
  OA22X1 U5037 ( .IN1(n5322), .IN2(n4171), .IN3(n6313), .IN4(n5332), .Q(n4170)
         );
  OA22X1 U5038 ( .IN1(n5965), .IN2(n5308), .IN3(n5315), .IN4(n4172), .Q(n4171)
         );
  OA22X1 U5039 ( .IN1(n5287), .IN2(n4173), .IN3(n6159), .IN4(n5298), .Q(n4172)
         );
  OA22X1 U5040 ( .IN1(n5950), .IN2(n5280), .IN3(n5283), .IN4(n6005), .Q(n4173)
         );
  OAI22X1 U5041 ( .IN1(n5341), .IN2(n4174), .IN3(n5981), .IN4(n5344), .QN(
        N10161) );
  OA22X1 U5042 ( .IN1(n5322), .IN2(n4175), .IN3(n6314), .IN4(n5332), .Q(n4174)
         );
  OA22X1 U5043 ( .IN1(n5966), .IN2(n5308), .IN3(n5312), .IN4(n4176), .Q(n4175)
         );
  OA22X1 U5044 ( .IN1(n5287), .IN2(n4177), .IN3(n6160), .IN4(n5298), .Q(n4176)
         );
  OA22X1 U5045 ( .IN1(n5951), .IN2(n5280), .IN3(n5283), .IN4(n6006), .Q(n4177)
         );
  OAI22X1 U5046 ( .IN1(n5341), .IN2(n4178), .IN3(n6375), .IN4(n5345), .QN(
        N10160) );
  OA22X1 U5047 ( .IN1(n5322), .IN2(n4179), .IN3(n6307), .IN4(n5332), .Q(n4178)
         );
  OA22X1 U5048 ( .IN1(n6221), .IN2(n5308), .IN3(n5315), .IN4(n4180), .Q(n4179)
         );
  OA22X1 U5049 ( .IN1(n5287), .IN2(n4181), .IN3(n6153), .IN4(n5298), .Q(n4180)
         );
  OA22X1 U5050 ( .IN1(n6067), .IN2(n5280), .IN3(n5283), .IN4(n5999), .Q(n4181)
         );
  OAI22X1 U5051 ( .IN1(n5341), .IN2(n4182), .IN3(n6372), .IN4(n5346), .QN(
        N10158) );
  OA22X1 U5052 ( .IN1(n5322), .IN2(n4183), .IN3(n6306), .IN4(n5332), .Q(n4182)
         );
  OA22X1 U5053 ( .IN1(n6218), .IN2(n5308), .IN3(n5310), .IN4(n4184), .Q(n4183)
         );
  OA22X1 U5054 ( .IN1(n5287), .IN2(n4185), .IN3(n6152), .IN4(n5298), .Q(n4184)
         );
  OA22X1 U5055 ( .IN1(n6064), .IN2(n5280), .IN3(n5283), .IN4(n5998), .Q(n4185)
         );
  OAI22X1 U5056 ( .IN1(n5341), .IN2(n4186), .IN3(n6377), .IN4(n5347), .QN(
        N10156) );
  OA22X1 U5057 ( .IN1(n5323), .IN2(n4187), .IN3(n6422), .IN4(n5332), .Q(n4186)
         );
  OA22X1 U5058 ( .IN1(n6223), .IN2(n5308), .IN3(n5311), .IN4(n4188), .Q(n4187)
         );
  OA22X1 U5059 ( .IN1(n5288), .IN2(n4189), .IN3(n6268), .IN4(n5298), .Q(n4188)
         );
  OA22X1 U5060 ( .IN1(n6069), .IN2(n5280), .IN3(n5283), .IN4(n6114), .Q(n4189)
         );
  OAI22X1 U5061 ( .IN1(n5341), .IN2(n4190), .IN3(n6378), .IN4(n5350), .QN(
        N10155) );
  OA22X1 U5062 ( .IN1(n5323), .IN2(n4191), .IN3(n6421), .IN4(n5332), .Q(n4190)
         );
  OA22X1 U5063 ( .IN1(n6224), .IN2(n5308), .IN3(n5313), .IN4(n4192), .Q(n4191)
         );
  OA22X1 U5064 ( .IN1(n5288), .IN2(n4193), .IN3(n6267), .IN4(n5298), .Q(n4192)
         );
  OA22X1 U5065 ( .IN1(n6070), .IN2(n5280), .IN3(n5283), .IN4(n6113), .Q(n4193)
         );
  OAI22X1 U5066 ( .IN1(n5341), .IN2(n4194), .IN3(n6379), .IN4(n5350), .QN(
        N10154) );
  OA22X1 U5067 ( .IN1(n5323), .IN2(n4195), .IN3(n6420), .IN4(n5332), .Q(n4194)
         );
  OA22X1 U5068 ( .IN1(n6225), .IN2(n5308), .IN3(n5311), .IN4(n4196), .Q(n4195)
         );
  OA22X1 U5069 ( .IN1(n5288), .IN2(n4197), .IN3(n6266), .IN4(n5298), .Q(n4196)
         );
  OA22X1 U5070 ( .IN1(n6071), .IN2(n5280), .IN3(n5283), .IN4(n6112), .Q(n4197)
         );
  OAI22X1 U5071 ( .IN1(n5341), .IN2(n4198), .IN3(n6380), .IN4(n5350), .QN(
        N10153) );
  OA22X1 U5072 ( .IN1(n5323), .IN2(n4199), .IN3(n6419), .IN4(n5332), .Q(n4198)
         );
  OA22X1 U5073 ( .IN1(n6226), .IN2(n5308), .IN3(n5311), .IN4(n4200), .Q(n4199)
         );
  OA22X1 U5074 ( .IN1(n5288), .IN2(n4201), .IN3(n6265), .IN4(n5298), .Q(n4200)
         );
  OA22X1 U5075 ( .IN1(n6072), .IN2(n5280), .IN3(n5283), .IN4(n6111), .Q(n4201)
         );
  OAI22X1 U5076 ( .IN1(n5341), .IN2(n4202), .IN3(n6381), .IN4(n5350), .QN(
        N10152) );
  OA22X1 U5077 ( .IN1(n5323), .IN2(n4203), .IN3(n6418), .IN4(n5332), .Q(n4202)
         );
  OA22X1 U5078 ( .IN1(n6227), .IN2(n5308), .IN3(n5311), .IN4(n4204), .Q(n4203)
         );
  OA22X1 U5079 ( .IN1(n5288), .IN2(n4205), .IN3(n6264), .IN4(n5298), .Q(n4204)
         );
  OA22X1 U5080 ( .IN1(n6073), .IN2(n5280), .IN3(n5282), .IN4(n6110), .Q(n4205)
         );
  OAI22X1 U5081 ( .IN1(n5341), .IN2(n4206), .IN3(n6382), .IN4(n5350), .QN(
        N10151) );
  OA22X1 U5082 ( .IN1(n5323), .IN2(n4207), .IN3(n6417), .IN4(n5332), .Q(n4206)
         );
  OA22X1 U5083 ( .IN1(n6228), .IN2(n5308), .IN3(n5311), .IN4(n4208), .Q(n4207)
         );
  OA22X1 U5084 ( .IN1(n5288), .IN2(n4209), .IN3(n6263), .IN4(n5298), .Q(n4208)
         );
  OA22X1 U5085 ( .IN1(n6074), .IN2(n5280), .IN3(n5199), .IN4(n6109), .Q(n4209)
         );
  OAI22X1 U5086 ( .IN1(n5341), .IN2(n4210), .IN3(n6383), .IN4(n5350), .QN(
        N10150) );
  OA22X1 U5087 ( .IN1(n5323), .IN2(n4211), .IN3(n6416), .IN4(n5332), .Q(n4210)
         );
  OA22X1 U5088 ( .IN1(n6229), .IN2(n5308), .IN3(n5311), .IN4(n4212), .Q(n4211)
         );
  OA22X1 U5089 ( .IN1(n5288), .IN2(n4213), .IN3(n6262), .IN4(n5298), .Q(n4212)
         );
  OA22X1 U5090 ( .IN1(n6075), .IN2(n5280), .IN3(n5199), .IN4(n6108), .Q(n4213)
         );
  OAI22X1 U5091 ( .IN1(n5341), .IN2(n4214), .IN3(n6385), .IN4(n5349), .QN(
        N10149) );
  OA22X1 U5092 ( .IN1(n5323), .IN2(n4215), .IN3(n6359), .IN4(n5332), .Q(n4214)
         );
  OA22X1 U5093 ( .IN1(n6231), .IN2(n5308), .IN3(n5312), .IN4(n4216), .Q(n4215)
         );
  OA22X1 U5094 ( .IN1(n5288), .IN2(n4217), .IN3(n6205), .IN4(n5298), .Q(n4216)
         );
  OA22X1 U5095 ( .IN1(n6077), .IN2(n5280), .IN3(n5199), .IN4(n6051), .Q(n4217)
         );
  OAI22X1 U5096 ( .IN1(n5341), .IN2(n4218), .IN3(n6386), .IN4(n5349), .QN(
        N10148) );
  OA22X1 U5097 ( .IN1(n5323), .IN2(n4219), .IN3(n6358), .IN4(n5333), .Q(n4218)
         );
  OA22X1 U5098 ( .IN1(n6232), .IN2(n5308), .IN3(n5312), .IN4(n4220), .Q(n4219)
         );
  OA22X1 U5099 ( .IN1(n5288), .IN2(n4221), .IN3(n6204), .IN4(n5298), .Q(n4220)
         );
  OA22X1 U5100 ( .IN1(n6078), .IN2(n5280), .IN3(n5199), .IN4(n6050), .Q(n4221)
         );
  OAI22X1 U5101 ( .IN1(n5341), .IN2(n4222), .IN3(n6387), .IN4(n5349), .QN(
        N10147) );
  OA22X1 U5102 ( .IN1(n5323), .IN2(n4223), .IN3(n6357), .IN4(n5333), .Q(n4222)
         );
  OA22X1 U5103 ( .IN1(n6233), .IN2(n5308), .IN3(n5312), .IN4(n4224), .Q(n4223)
         );
  OA22X1 U5104 ( .IN1(n5288), .IN2(n4225), .IN3(n6203), .IN4(n5303), .Q(n4224)
         );
  OA22X1 U5105 ( .IN1(n6079), .IN2(n5280), .IN3(n5199), .IN4(n6049), .Q(n4225)
         );
  OAI22X1 U5106 ( .IN1(n5341), .IN2(n4226), .IN3(n6388), .IN4(n5349), .QN(
        N10146) );
  OA22X1 U5107 ( .IN1(n5323), .IN2(n4227), .IN3(n6356), .IN4(n5333), .Q(n4226)
         );
  OA22X1 U5108 ( .IN1(n6234), .IN2(n5308), .IN3(n5312), .IN4(n4228), .Q(n4227)
         );
  OA22X1 U5109 ( .IN1(n5288), .IN2(n4229), .IN3(n6202), .IN4(n5284), .Q(n4228)
         );
  OA22X1 U5110 ( .IN1(n6080), .IN2(n5280), .IN3(n5199), .IN4(n6048), .Q(n4229)
         );
  OAI22X1 U5111 ( .IN1(n5341), .IN2(n4230), .IN3(n6389), .IN4(n5349), .QN(
        N10145) );
  OA22X1 U5112 ( .IN1(n5323), .IN2(n4231), .IN3(n6355), .IN4(n5333), .Q(n4230)
         );
  OA22X1 U5113 ( .IN1(n6235), .IN2(n5308), .IN3(n5312), .IN4(n4232), .Q(n4231)
         );
  OA22X1 U5114 ( .IN1(n5288), .IN2(n4233), .IN3(n6201), .IN4(n5285), .Q(n4232)
         );
  OA22X1 U5115 ( .IN1(n6081), .IN2(n5280), .IN3(n5282), .IN4(n6047), .Q(n4233)
         );
  OAI22X1 U5116 ( .IN1(n5341), .IN2(n4234), .IN3(n6390), .IN4(n5349), .QN(
        N10144) );
  OA22X1 U5117 ( .IN1(n5324), .IN2(n4235), .IN3(n6354), .IN4(n5333), .Q(n4234)
         );
  OA22X1 U5118 ( .IN1(n6236), .IN2(n5308), .IN3(n5313), .IN4(n4236), .Q(n4235)
         );
  OA22X1 U5119 ( .IN1(n5289), .IN2(n4237), .IN3(n6200), .IN4(n5284), .Q(n4236)
         );
  OA22X1 U5120 ( .IN1(n6082), .IN2(n5280), .IN3(n5199), .IN4(n6046), .Q(n4237)
         );
  OAI22X1 U5121 ( .IN1(n5341), .IN2(n4238), .IN3(n6391), .IN4(n5346), .QN(
        N10143) );
  OA22X1 U5122 ( .IN1(n5324), .IN2(n4239), .IN3(n6353), .IN4(n5333), .Q(n4238)
         );
  OA22X1 U5123 ( .IN1(n6237), .IN2(n5308), .IN3(n5313), .IN4(n4240), .Q(n4239)
         );
  OA22X1 U5124 ( .IN1(n5289), .IN2(n4241), .IN3(n6199), .IN4(n5285), .Q(n4240)
         );
  OA22X1 U5125 ( .IN1(n6083), .IN2(n5280), .IN3(n5199), .IN4(n6045), .Q(n4241)
         );
  OAI22X1 U5126 ( .IN1(n5341), .IN2(n4242), .IN3(n6400), .IN4(n5347), .QN(
        N10142) );
  OA22X1 U5127 ( .IN1(n5324), .IN2(n4243), .IN3(n6415), .IN4(n5333), .Q(n4242)
         );
  OA22X1 U5128 ( .IN1(n6246), .IN2(n5308), .IN3(n5313), .IN4(n4244), .Q(n4243)
         );
  OA22X1 U5129 ( .IN1(n5289), .IN2(n4245), .IN3(n6261), .IN4(n5284), .Q(n4244)
         );
  OA22X1 U5130 ( .IN1(n6092), .IN2(n5280), .IN3(n5199), .IN4(n6107), .Q(n4245)
         );
  OAI22X1 U5131 ( .IN1(n5341), .IN2(n4246), .IN3(n6406), .IN4(n5343), .QN(
        N10141) );
  OA22X1 U5132 ( .IN1(n5324), .IN2(n4247), .IN3(n6414), .IN4(n5333), .Q(n4246)
         );
  OA22X1 U5133 ( .IN1(n6252), .IN2(n5308), .IN3(n5313), .IN4(n4248), .Q(n4247)
         );
  OA22X1 U5134 ( .IN1(n5289), .IN2(n4249), .IN3(n6260), .IN4(n5285), .Q(n4248)
         );
  OA22X1 U5135 ( .IN1(n6098), .IN2(n5280), .IN3(n5199), .IN4(n6106), .Q(n4249)
         );
  OAI22X1 U5136 ( .IN1(n5341), .IN2(n4250), .IN3(n6407), .IN4(n5348), .QN(
        N10140) );
  OA22X1 U5137 ( .IN1(n5324), .IN2(n4251), .IN3(n6413), .IN4(n5333), .Q(n4250)
         );
  OA22X1 U5138 ( .IN1(n6253), .IN2(n5308), .IN3(n5313), .IN4(n4252), .Q(n4251)
         );
  OA22X1 U5139 ( .IN1(n5289), .IN2(n4253), .IN3(n6259), .IN4(n5284), .Q(n4252)
         );
  OA22X1 U5140 ( .IN1(n6099), .IN2(n5280), .IN3(n5199), .IN4(n6105), .Q(n4253)
         );
  OAI22X1 U5141 ( .IN1(n5341), .IN2(n4254), .IN3(n6408), .IN4(n5349), .QN(
        N10139) );
  OA22X1 U5142 ( .IN1(n5324), .IN2(n4255), .IN3(n6412), .IN4(n5333), .Q(n4254)
         );
  OA22X1 U5143 ( .IN1(n6254), .IN2(n5308), .IN3(n5317), .IN4(n4256), .Q(n4255)
         );
  OA22X1 U5144 ( .IN1(n5289), .IN2(n4257), .IN3(n6258), .IN4(n5285), .Q(n4256)
         );
  OA22X1 U5145 ( .IN1(n6100), .IN2(n5280), .IN3(n5199), .IN4(n6104), .Q(n4257)
         );
  OAI22X1 U5146 ( .IN1(n5341), .IN2(n4258), .IN3(n6409), .IN4(n5350), .QN(
        N10138) );
  OA22X1 U5147 ( .IN1(n5324), .IN2(n4259), .IN3(n6411), .IN4(n5333), .Q(n4258)
         );
  OA22X1 U5148 ( .IN1(n6255), .IN2(n5308), .IN3(n5312), .IN4(n4260), .Q(n4259)
         );
  OA22X1 U5149 ( .IN1(n5289), .IN2(n4261), .IN3(n6257), .IN4(n5284), .Q(n4260)
         );
  OA22X1 U5150 ( .IN1(n6101), .IN2(n5280), .IN3(n5199), .IN4(n6103), .Q(n4261)
         );
  OAI22X1 U5151 ( .IN1(n5341), .IN2(n4262), .IN3(n6401), .IN4(n5348), .QN(
        N10137) );
  OA22X1 U5152 ( .IN1(n5324), .IN2(n4263), .IN3(n6410), .IN4(n5333), .Q(n4262)
         );
  OA22X1 U5153 ( .IN1(n6247), .IN2(n5308), .IN3(n5316), .IN4(n4264), .Q(n4263)
         );
  OA22X1 U5154 ( .IN1(n5289), .IN2(n4265), .IN3(n6256), .IN4(n5285), .Q(n4264)
         );
  OA22X1 U5155 ( .IN1(n6093), .IN2(n5280), .IN3(n5199), .IN4(n6102), .Q(n4265)
         );
  OAI22X1 U5156 ( .IN1(n5341), .IN2(n4266), .IN3(n6399), .IN4(n5348), .QN(
        N10136) );
  OA22X1 U5157 ( .IN1(n5324), .IN2(n4267), .IN3(n6352), .IN4(n5333), .Q(n4266)
         );
  OA22X1 U5158 ( .IN1(n6244), .IN2(n5308), .IN3(n5315), .IN4(n4268), .Q(n4267)
         );
  OA22X1 U5159 ( .IN1(n5289), .IN2(n4269), .IN3(n6198), .IN4(n5284), .Q(n4268)
         );
  OA22X1 U5160 ( .IN1(n6090), .IN2(n5280), .IN3(n5199), .IN4(n6044), .Q(n4269)
         );
  OAI22X1 U5161 ( .IN1(n5341), .IN2(n4270), .IN3(n6398), .IN4(n5348), .QN(
        N10135) );
  OA22X1 U5162 ( .IN1(n5324), .IN2(n4271), .IN3(n6402), .IN4(n5333), .Q(n4270)
         );
  OA22X1 U5163 ( .IN1(n6243), .IN2(n5308), .IN3(n5313), .IN4(n4272), .Q(n4271)
         );
  OA22X1 U5164 ( .IN1(n5289), .IN2(n4273), .IN3(n6248), .IN4(n5285), .Q(n4272)
         );
  OA22X1 U5165 ( .IN1(n6089), .IN2(n5280), .IN3(n5199), .IN4(n6094), .Q(n4273)
         );
  OAI22X1 U5166 ( .IN1(n5342), .IN2(n4274), .IN3(n6397), .IN4(n5348), .QN(
        N10134) );
  OA22X1 U5167 ( .IN1(n5324), .IN2(n4275), .IN3(n6403), .IN4(n5333), .Q(n4274)
         );
  OA22X1 U5168 ( .IN1(n6242), .IN2(n5308), .IN3(n5311), .IN4(n4276), .Q(n4275)
         );
  OA22X1 U5169 ( .IN1(n5289), .IN2(n4277), .IN3(n6249), .IN4(n5284), .Q(n4276)
         );
  OA22X1 U5170 ( .IN1(n6091), .IN2(n5280), .IN3(n5199), .IN4(n6095), .Q(n4277)
         );
  OAI22X1 U5171 ( .IN1(n5342), .IN2(n4278), .IN3(n6396), .IN4(n5348), .QN(
        N10133) );
  OA22X1 U5172 ( .IN1(n5324), .IN2(n4279), .IN3(n6404), .IN4(n5334), .Q(n4278)
         );
  OA22X1 U5173 ( .IN1(n6241), .IN2(n5308), .IN3(n5315), .IN4(n4280), .Q(n4279)
         );
  OA22X1 U5174 ( .IN1(n5289), .IN2(n4281), .IN3(n6250), .IN4(n5284), .Q(n4280)
         );
  OA22X1 U5175 ( .IN1(n6088), .IN2(n5280), .IN3(n5199), .IN4(n6096), .Q(n4281)
         );
  OAI22X1 U5176 ( .IN1(n5342), .IN2(n4282), .IN3(n6398), .IN4(n5348), .QN(
        N10132) );
  OA22X1 U5177 ( .IN1(n5325), .IN2(n4283), .IN3(n6405), .IN4(n5334), .Q(n4282)
         );
  OA22X1 U5178 ( .IN1(n6245), .IN2(n5308), .IN3(n5310), .IN4(n4284), .Q(n4283)
         );
  OA22X1 U5179 ( .IN1(n5290), .IN2(n4285), .IN3(n6251), .IN4(n5299), .Q(n4284)
         );
  OA22X1 U5180 ( .IN1(n6087), .IN2(n5280), .IN3(n5199), .IN4(n6097), .Q(n4285)
         );
  OAI22X1 U5181 ( .IN1(n5342), .IN2(n4286), .IN3(n6394), .IN4(n5347), .QN(
        N10131) );
  OA22X1 U5182 ( .IN1(n5325), .IN2(n4287), .IN3(n6393), .IN4(n5334), .Q(n4286)
         );
  OA22X1 U5183 ( .IN1(n6240), .IN2(n5308), .IN3(n5311), .IN4(n4288), .Q(n4287)
         );
  OA22X1 U5184 ( .IN1(n5290), .IN2(n4289), .IN3(n6239), .IN4(n5299), .Q(n4288)
         );
  OA22X1 U5185 ( .IN1(n6086), .IN2(n5280), .IN3(n5199), .IN4(n6085), .Q(n4289)
         );
  OAI22X1 U5186 ( .IN1(n5342), .IN2(n4290), .IN3(n6361), .IN4(n5347), .QN(
        N10130) );
  OA22X1 U5187 ( .IN1(n5325), .IN2(n4291), .IN3(n6360), .IN4(n5334), .Q(n4290)
         );
  OA22X1 U5188 ( .IN1(n6207), .IN2(n5308), .IN3(n5313), .IN4(n4292), .Q(n4291)
         );
  OA22X1 U5189 ( .IN1(n5290), .IN2(n4293), .IN3(n6206), .IN4(n5299), .Q(n4292)
         );
  OA22X1 U5190 ( .IN1(n6053), .IN2(n5280), .IN3(n5199), .IN4(n6052), .Q(n4293)
         );
  OAI22X1 U5191 ( .IN1(n5342), .IN2(n4294), .IN3(n6350), .IN4(n5347), .QN(
        N10129) );
  OA22X1 U5192 ( .IN1(n5325), .IN2(n4295), .IN3(n6351), .IN4(n5334), .Q(n4294)
         );
  OA22X1 U5193 ( .IN1(n6196), .IN2(n5308), .IN3(n5314), .IN4(n4296), .Q(n4295)
         );
  OA22X1 U5194 ( .IN1(n5290), .IN2(n4297), .IN3(n6197), .IN4(n5299), .Q(n4296)
         );
  OA22X1 U5195 ( .IN1(n6042), .IN2(n5279), .IN3(n5199), .IN4(n6043), .Q(n4297)
         );
  OAI22X1 U5196 ( .IN1(n5342), .IN2(n4298), .IN3(n6395), .IN4(n5347), .QN(
        N10128) );
  OA22X1 U5197 ( .IN1(n5325), .IN2(n4299), .IN3(n6392), .IN4(n5334), .Q(n4298)
         );
  OA22X1 U5198 ( .IN1(n6244), .IN2(n5307), .IN3(n5314), .IN4(n4300), .Q(n4299)
         );
  OA22X1 U5199 ( .IN1(n5290), .IN2(n4301), .IN3(n6238), .IN4(n5299), .Q(n4300)
         );
  OA22X1 U5200 ( .IN1(n6090), .IN2(n5279), .IN3(n5199), .IN4(n6084), .Q(n4301)
         );
  OAI22X1 U5201 ( .IN1(n5342), .IN2(n4302), .IN3(n6423), .IN4(n5347), .QN(
        N10127) );
  OA22X1 U5202 ( .IN1(n5325), .IN2(n4303), .IN3(n6423), .IN4(n5334), .Q(n4302)
         );
  OA22X1 U5203 ( .IN1(n6269), .IN2(n5307), .IN3(n5314), .IN4(n4304), .Q(n4303)
         );
  OA22X1 U5204 ( .IN1(n5290), .IN2(n4305), .IN3(n6269), .IN4(n5299), .Q(n4304)
         );
  OA22X1 U5205 ( .IN1(n6115), .IN2(n5279), .IN3(n5199), .IN4(n6115), .Q(n4305)
         );
  OAI22X1 U5206 ( .IN1(n5342), .IN2(n4306), .IN3(n6424), .IN4(n5347), .QN(
        N10126) );
  OA22X1 U5207 ( .IN1(n5325), .IN2(n4307), .IN3(n6424), .IN4(n5334), .Q(n4306)
         );
  OA22X1 U5208 ( .IN1(n6270), .IN2(n5307), .IN3(n5314), .IN4(n4308), .Q(n4307)
         );
  OA22X1 U5209 ( .IN1(n5290), .IN2(n4309), .IN3(n6270), .IN4(n5299), .Q(n4308)
         );
  OA22X1 U5210 ( .IN1(n6116), .IN2(n5279), .IN3(n5199), .IN4(n6116), .Q(n4309)
         );
  OAI22X1 U5211 ( .IN1(n5342), .IN2(n4310), .IN3(n6425), .IN4(n5346), .QN(
        N10125) );
  OA22X1 U5212 ( .IN1(n5325), .IN2(n4311), .IN3(n6425), .IN4(n5334), .Q(n4310)
         );
  OA22X1 U5213 ( .IN1(n6271), .IN2(n5307), .IN3(n5314), .IN4(n4312), .Q(n4311)
         );
  OA22X1 U5214 ( .IN1(n5290), .IN2(n4313), .IN3(n6271), .IN4(n5299), .Q(n4312)
         );
  OA22X1 U5215 ( .IN1(n6117), .IN2(n5279), .IN3(n5199), .IN4(n6117), .Q(n4313)
         );
  OAI22X1 U5216 ( .IN1(n5342), .IN2(n4314), .IN3(n6426), .IN4(n5346), .QN(
        N10124) );
  OA22X1 U5217 ( .IN1(n5325), .IN2(n4315), .IN3(n6426), .IN4(n5334), .Q(n4314)
         );
  OA22X1 U5218 ( .IN1(n6272), .IN2(n5307), .IN3(n5315), .IN4(n4316), .Q(n4315)
         );
  OA22X1 U5219 ( .IN1(n5290), .IN2(n4317), .IN3(n6272), .IN4(n5299), .Q(n4316)
         );
  OA22X1 U5220 ( .IN1(n6118), .IN2(n5279), .IN3(n5199), .IN4(n6118), .Q(n4317)
         );
  OAI22X1 U5221 ( .IN1(n5342), .IN2(n4318), .IN3(n6427), .IN4(n5346), .QN(
        N10123) );
  OA22X1 U5222 ( .IN1(n5325), .IN2(n4319), .IN3(n6427), .IN4(n5334), .Q(n4318)
         );
  OA22X1 U5223 ( .IN1(n6273), .IN2(n5307), .IN3(n5313), .IN4(n4320), .Q(n4319)
         );
  OA22X1 U5224 ( .IN1(n5290), .IN2(n4321), .IN3(n6273), .IN4(n5299), .Q(n4320)
         );
  OA22X1 U5225 ( .IN1(n6119), .IN2(n5279), .IN3(n5199), .IN4(n6119), .Q(n4321)
         );
  OAI22X1 U5226 ( .IN1(n5342), .IN2(n4322), .IN3(n6428), .IN4(n5346), .QN(
        N10122) );
  OA22X1 U5227 ( .IN1(n5325), .IN2(n4323), .IN3(n6428), .IN4(n5334), .Q(n4322)
         );
  OA22X1 U5228 ( .IN1(n6274), .IN2(n5307), .IN3(n5316), .IN4(n4324), .Q(n4323)
         );
  OA22X1 U5229 ( .IN1(n5290), .IN2(n4325), .IN3(n6274), .IN4(n5299), .Q(n4324)
         );
  OA22X1 U5230 ( .IN1(n6120), .IN2(n5279), .IN3(n5199), .IN4(n6120), .Q(n4325)
         );
  OAI22X1 U5231 ( .IN1(n5342), .IN2(n4326), .IN3(n6429), .IN4(n5346), .QN(
        N10121) );
  OA22X1 U5232 ( .IN1(n5325), .IN2(n4327), .IN3(n6429), .IN4(n5334), .Q(n4326)
         );
  OA22X1 U5233 ( .IN1(n6275), .IN2(n5307), .IN3(n5316), .IN4(n4328), .Q(n4327)
         );
  OA22X1 U5234 ( .IN1(n5290), .IN2(n4329), .IN3(n6275), .IN4(n5299), .Q(n4328)
         );
  OA22X1 U5235 ( .IN1(n6121), .IN2(n5279), .IN3(n5199), .IN4(n6121), .Q(n4329)
         );
  OAI22X1 U5236 ( .IN1(n5342), .IN2(n4330), .IN3(n6430), .IN4(n5346), .QN(
        N10120) );
  OA22X1 U5237 ( .IN1(n5326), .IN2(n4331), .IN3(n6430), .IN4(n5334), .Q(n4330)
         );
  OA22X1 U5238 ( .IN1(n6276), .IN2(n5307), .IN3(n5314), .IN4(n4332), .Q(n4331)
         );
  OA22X1 U5239 ( .IN1(n5291), .IN2(n4333), .IN3(n6276), .IN4(n5299), .Q(n4332)
         );
  OA22X1 U5240 ( .IN1(n6122), .IN2(n5279), .IN3(n5199), .IN4(n6122), .Q(n4333)
         );
  OAI22X1 U5241 ( .IN1(n5342), .IN2(n4334), .IN3(n6431), .IN4(n5345), .QN(
        N10119) );
  OA22X1 U5242 ( .IN1(n5326), .IN2(n4335), .IN3(n6431), .IN4(n5335), .Q(n4334)
         );
  OA22X1 U5243 ( .IN1(n6277), .IN2(n5307), .IN3(n5315), .IN4(n4336), .Q(n4335)
         );
  OA22X1 U5244 ( .IN1(n5291), .IN2(n4337), .IN3(n6277), .IN4(n5299), .Q(n4336)
         );
  OA22X1 U5245 ( .IN1(n6123), .IN2(n5279), .IN3(n5282), .IN4(n6123), .Q(n4337)
         );
  OAI22X1 U5246 ( .IN1(n5342), .IN2(n4338), .IN3(n6432), .IN4(n5345), .QN(
        N10118) );
  OA22X1 U5247 ( .IN1(n5326), .IN2(n4339), .IN3(n6432), .IN4(n5335), .Q(n4338)
         );
  OA22X1 U5248 ( .IN1(n6278), .IN2(n5307), .IN3(n5315), .IN4(n4340), .Q(n4339)
         );
  OA22X1 U5249 ( .IN1(n5291), .IN2(n4341), .IN3(n6278), .IN4(n5300), .Q(n4340)
         );
  OA22X1 U5250 ( .IN1(n6124), .IN2(n5279), .IN3(n5282), .IN4(n6124), .Q(n4341)
         );
  OAI22X1 U5251 ( .IN1(n5342), .IN2(n4342), .IN3(n6433), .IN4(n5345), .QN(
        N10117) );
  OA22X1 U5252 ( .IN1(n5326), .IN2(n4343), .IN3(n6433), .IN4(n5335), .Q(n4342)
         );
  OA22X1 U5253 ( .IN1(n6279), .IN2(n5307), .IN3(n5315), .IN4(n4344), .Q(n4343)
         );
  OA22X1 U5254 ( .IN1(n5291), .IN2(n4345), .IN3(n6279), .IN4(n5300), .Q(n4344)
         );
  OA22X1 U5255 ( .IN1(n6125), .IN2(n5279), .IN3(n5282), .IN4(n6125), .Q(n4345)
         );
  OAI22X1 U5256 ( .IN1(n5342), .IN2(n4346), .IN3(n6434), .IN4(n5345), .QN(
        N10116) );
  OA22X1 U5257 ( .IN1(n5326), .IN2(n4347), .IN3(n6434), .IN4(n5335), .Q(n4346)
         );
  OA22X1 U5258 ( .IN1(n6280), .IN2(n5307), .IN3(n5315), .IN4(n4348), .Q(n4347)
         );
  OA22X1 U5259 ( .IN1(n5291), .IN2(n4349), .IN3(n6280), .IN4(n5300), .Q(n4348)
         );
  OA22X1 U5260 ( .IN1(n6126), .IN2(n5279), .IN3(n5282), .IN4(n6126), .Q(n4349)
         );
  OAI22X1 U5261 ( .IN1(n5342), .IN2(n4350), .IN3(n6435), .IN4(n5345), .QN(
        N10115) );
  OA22X1 U5262 ( .IN1(n5326), .IN2(n4351), .IN3(n6435), .IN4(n5335), .Q(n4350)
         );
  OA22X1 U5263 ( .IN1(n6281), .IN2(n5307), .IN3(n5315), .IN4(n4352), .Q(n4351)
         );
  OA22X1 U5264 ( .IN1(n5291), .IN2(n4353), .IN3(n6281), .IN4(n5300), .Q(n4352)
         );
  OA22X1 U5265 ( .IN1(n6127), .IN2(n5279), .IN3(n5282), .IN4(n6127), .Q(n4353)
         );
  OAI22X1 U5266 ( .IN1(n5342), .IN2(n4354), .IN3(n6436), .IN4(n5345), .QN(
        N10114) );
  OA22X1 U5267 ( .IN1(n5326), .IN2(n4355), .IN3(n6436), .IN4(n5335), .Q(n4354)
         );
  OA22X1 U5268 ( .IN1(n6282), .IN2(n5307), .IN3(n5316), .IN4(n4356), .Q(n4355)
         );
  OA22X1 U5269 ( .IN1(n5291), .IN2(n4357), .IN3(n6282), .IN4(n5300), .Q(n4356)
         );
  OA22X1 U5270 ( .IN1(n6128), .IN2(n5279), .IN3(n5282), .IN4(n6128), .Q(n4357)
         );
  OAI22X1 U5271 ( .IN1(n5342), .IN2(n4358), .IN3(n6437), .IN4(n5344), .QN(
        N10113) );
  OA22X1 U5272 ( .IN1(n5326), .IN2(n4359), .IN3(n6437), .IN4(n5335), .Q(n4358)
         );
  OA22X1 U5273 ( .IN1(n6283), .IN2(n5307), .IN3(n5316), .IN4(n4360), .Q(n4359)
         );
  OA22X1 U5274 ( .IN1(n5291), .IN2(n4361), .IN3(n6283), .IN4(n5300), .Q(n4360)
         );
  OA22X1 U5275 ( .IN1(n6129), .IN2(n5279), .IN3(n5282), .IN4(n6129), .Q(n4361)
         );
  OAI22X1 U5276 ( .IN1(n5342), .IN2(n4362), .IN3(n6438), .IN4(n5344), .QN(
        N10112) );
  OA22X1 U5277 ( .IN1(n5326), .IN2(n4363), .IN3(n6438), .IN4(n5335), .Q(n4362)
         );
  OA22X1 U5278 ( .IN1(n6284), .IN2(n5307), .IN3(n5316), .IN4(n4364), .Q(n4363)
         );
  OA22X1 U5279 ( .IN1(n5291), .IN2(n4365), .IN3(n6284), .IN4(n5300), .Q(n4364)
         );
  OA22X1 U5280 ( .IN1(n6130), .IN2(n5279), .IN3(n5282), .IN4(n6130), .Q(n4365)
         );
  OAI22X1 U5281 ( .IN1(n5342), .IN2(n4366), .IN3(n6439), .IN4(n5344), .QN(
        N10111) );
  OA22X1 U5282 ( .IN1(n5326), .IN2(n4367), .IN3(n6439), .IN4(n5335), .Q(n4366)
         );
  OA22X1 U5283 ( .IN1(n6285), .IN2(n5307), .IN3(n5316), .IN4(n4368), .Q(n4367)
         );
  OA22X1 U5284 ( .IN1(n5291), .IN2(n4369), .IN3(n6285), .IN4(n5300), .Q(n4368)
         );
  OA22X1 U5285 ( .IN1(n6131), .IN2(n5279), .IN3(n5282), .IN4(n6131), .Q(n4369)
         );
  OAI22X1 U5286 ( .IN1(n5342), .IN2(n4370), .IN3(n6440), .IN4(n5344), .QN(
        N10110) );
  OA22X1 U5287 ( .IN1(n5326), .IN2(n4371), .IN3(n6440), .IN4(n5335), .Q(n4370)
         );
  OA22X1 U5288 ( .IN1(n6286), .IN2(n5307), .IN3(n5316), .IN4(n4372), .Q(n4371)
         );
  OA22X1 U5289 ( .IN1(n5291), .IN2(n4373), .IN3(n6286), .IN4(n5300), .Q(n4372)
         );
  OA22X1 U5290 ( .IN1(n6132), .IN2(n5279), .IN3(n5282), .IN4(n6132), .Q(n4373)
         );
  OAI22X1 U5291 ( .IN1(n5342), .IN2(n4374), .IN3(n6441), .IN4(n5344), .QN(
        N10109) );
  OA22X1 U5292 ( .IN1(n5326), .IN2(n4375), .IN3(n6441), .IN4(n5335), .Q(n4374)
         );
  OA22X1 U5293 ( .IN1(n6287), .IN2(n5307), .IN3(n5317), .IN4(n4376), .Q(n4375)
         );
  OA22X1 U5294 ( .IN1(n5291), .IN2(n4377), .IN3(n6287), .IN4(n5300), .Q(n4376)
         );
  OA22X1 U5295 ( .IN1(n6133), .IN2(n5279), .IN3(n5282), .IN4(n6133), .Q(n4377)
         );
  OAI22X1 U5296 ( .IN1(n5342), .IN2(n4378), .IN3(n6442), .IN4(n5344), .QN(
        N10108) );
  OA22X1 U5297 ( .IN1(n5327), .IN2(n4379), .IN3(n6442), .IN4(n5335), .Q(n4378)
         );
  OA22X1 U5298 ( .IN1(n6288), .IN2(n5307), .IN3(n5313), .IN4(n4380), .Q(n4379)
         );
  OA22X1 U5299 ( .IN1(n5292), .IN2(n4381), .IN3(n6288), .IN4(n5300), .Q(n4380)
         );
  OA22X1 U5300 ( .IN1(n6134), .IN2(n5279), .IN3(n5282), .IN4(n6134), .Q(n4381)
         );
  OAI22X1 U5301 ( .IN1(n5342), .IN2(n4382), .IN3(n6443), .IN4(n5345), .QN(
        N10106) );
  OA22X1 U5302 ( .IN1(n5327), .IN2(n4383), .IN3(n6443), .IN4(n5335), .Q(n4382)
         );
  OA22X1 U5303 ( .IN1(n6289), .IN2(n5307), .IN3(n5316), .IN4(n4384), .Q(n4383)
         );
  OA22X1 U5304 ( .IN1(n5292), .IN2(n4385), .IN3(n6289), .IN4(n5300), .Q(n4384)
         );
  OA22X1 U5305 ( .IN1(n6135), .IN2(n5279), .IN3(n5282), .IN4(n6135), .Q(n4385)
         );
  OAI22X1 U5306 ( .IN1(n5342), .IN2(n4386), .IN3(n6444), .IN4(n5344), .QN(
        N10105) );
  OA22X1 U5307 ( .IN1(n5327), .IN2(n4387), .IN3(n6444), .IN4(n5335), .Q(n4386)
         );
  OA22X1 U5308 ( .IN1(n6290), .IN2(n5307), .IN3(n5312), .IN4(n4388), .Q(n4387)
         );
  OA22X1 U5309 ( .IN1(n5292), .IN2(n4389), .IN3(n6290), .IN4(n5300), .Q(n4388)
         );
  OA22X1 U5310 ( .IN1(n6136), .IN2(n5279), .IN3(n5282), .IN4(n6136), .Q(n4389)
         );
  OAI22X1 U5311 ( .IN1(n5342), .IN2(n4390), .IN3(n6445), .IN4(n5346), .QN(
        N10104) );
  OA22X1 U5312 ( .IN1(n5327), .IN2(n4391), .IN3(n6445), .IN4(n5335), .Q(n4390)
         );
  OA22X1 U5313 ( .IN1(n6291), .IN2(n5307), .IN3(n5317), .IN4(n4392), .Q(n4391)
         );
  OA22X1 U5314 ( .IN1(n5292), .IN2(n4393), .IN3(n6291), .IN4(n5300), .Q(n4392)
         );
  OA22X1 U5315 ( .IN1(n6137), .IN2(n5279), .IN3(n5282), .IN4(n6137), .Q(n4393)
         );
  OAI22X1 U5316 ( .IN1(n5342), .IN2(n4394), .IN3(n6446), .IN4(n5347), .QN(
        N10103) );
  OA22X1 U5317 ( .IN1(n5327), .IN2(n4395), .IN3(n6446), .IN4(n5336), .Q(n4394)
         );
  OA22X1 U5318 ( .IN1(n6292), .IN2(n5307), .IN3(n5315), .IN4(n4396), .Q(n4395)
         );
  OA22X1 U5319 ( .IN1(n5292), .IN2(n4397), .IN3(n6292), .IN4(n5300), .Q(n4396)
         );
  OA22X1 U5320 ( .IN1(n6138), .IN2(n5279), .IN3(n5282), .IN4(n6138), .Q(n4397)
         );
  OAI22X1 U5321 ( .IN1(n5342), .IN2(n4398), .IN3(n6447), .IN4(n5343), .QN(
        N10102) );
  OA22X1 U5322 ( .IN1(n5327), .IN2(n4399), .IN3(n6447), .IN4(n5336), .Q(n4398)
         );
  OA22X1 U5323 ( .IN1(n6293), .IN2(n5307), .IN3(n5310), .IN4(n4400), .Q(n4399)
         );
  OA22X1 U5324 ( .IN1(n5292), .IN2(n4401), .IN3(n6293), .IN4(n5301), .Q(n4400)
         );
  OA22X1 U5325 ( .IN1(n6139), .IN2(n5279), .IN3(n5282), .IN4(n6139), .Q(n4401)
         );
  OAI22X1 U5326 ( .IN1(n5342), .IN2(n4402), .IN3(n6448), .IN4(n5348), .QN(
        N10101) );
  OA22X1 U5327 ( .IN1(n5327), .IN2(n4403), .IN3(n6448), .IN4(n5336), .Q(n4402)
         );
  OA22X1 U5328 ( .IN1(n6294), .IN2(n5307), .IN3(n5311), .IN4(n4404), .Q(n4403)
         );
  OA22X1 U5329 ( .IN1(n5292), .IN2(n4405), .IN3(n6294), .IN4(n5301), .Q(n4404)
         );
  OA22X1 U5330 ( .IN1(n6140), .IN2(n5279), .IN3(n5282), .IN4(n6140), .Q(n4405)
         );
  OAI22X1 U5331 ( .IN1(n5342), .IN2(n4406), .IN3(n6449), .IN4(n5343), .QN(
        N10100) );
  OA22X1 U5332 ( .IN1(n5327), .IN2(n4407), .IN3(n6449), .IN4(n5336), .Q(n4406)
         );
  OA22X1 U5333 ( .IN1(n6295), .IN2(n5307), .IN3(n5313), .IN4(n4408), .Q(n4407)
         );
  OA22X1 U5334 ( .IN1(n5292), .IN2(n4409), .IN3(n6295), .IN4(n5301), .Q(n4408)
         );
  OA22X1 U5335 ( .IN1(n6141), .IN2(n5279), .IN3(n5282), .IN4(n6141), .Q(n4409)
         );
  OAI22X1 U5336 ( .IN1(n5342), .IN2(n4410), .IN3(n6450), .IN4(n5343), .QN(
        N10099) );
  OA22X1 U5337 ( .IN1(n5327), .IN2(n4411), .IN3(n6450), .IN4(n5336), .Q(n4410)
         );
  OA22X1 U5338 ( .IN1(n6296), .IN2(n5307), .IN3(n5316), .IN4(n4412), .Q(n4411)
         );
  OA22X1 U5339 ( .IN1(n5292), .IN2(n4413), .IN3(n6296), .IN4(n5301), .Q(n4412)
         );
  OA22X1 U5340 ( .IN1(n6142), .IN2(n5279), .IN3(n5282), .IN4(n6142), .Q(n4413)
         );
  OAI22X1 U5341 ( .IN1(n5342), .IN2(n4414), .IN3(n6451), .IN4(n5343), .QN(
        N10098) );
  OA22X1 U5342 ( .IN1(n5327), .IN2(n4415), .IN3(n6451), .IN4(n5336), .Q(n4414)
         );
  OA22X1 U5343 ( .IN1(n6297), .IN2(n5307), .IN3(n5317), .IN4(n4416), .Q(n4415)
         );
  OA22X1 U5344 ( .IN1(n5292), .IN2(n4417), .IN3(n6297), .IN4(n5301), .Q(n4416)
         );
  OA22X1 U5345 ( .IN1(n6143), .IN2(n5279), .IN3(n5282), .IN4(n6143), .Q(n4417)
         );
  OAI22X1 U5346 ( .IN1(n5342), .IN2(n4418), .IN3(n6452), .IN4(n5343), .QN(
        N10097) );
  OA22X1 U5347 ( .IN1(n5327), .IN2(n4419), .IN3(n6452), .IN4(n5336), .Q(n4418)
         );
  OA22X1 U5348 ( .IN1(n6298), .IN2(n5307), .IN3(n5317), .IN4(n4420), .Q(n4419)
         );
  OA22X1 U5349 ( .IN1(n5292), .IN2(n4421), .IN3(n6298), .IN4(n5301), .Q(n4420)
         );
  OA22X1 U5350 ( .IN1(n6144), .IN2(n5279), .IN3(n5282), .IN4(n6144), .Q(n4421)
         );
  OAI22X1 U5351 ( .IN1(n5342), .IN2(n4422), .IN3(n6453), .IN4(n5343), .QN(
        N10096) );
  OA22X1 U5352 ( .IN1(n5327), .IN2(n4423), .IN3(n6453), .IN4(n5336), .Q(n4422)
         );
  OA22X1 U5353 ( .IN1(n6299), .IN2(n5307), .IN3(n5317), .IN4(n4424), .Q(n4423)
         );
  OA22X1 U5354 ( .IN1(n5292), .IN2(n4425), .IN3(n6299), .IN4(n5301), .Q(n4424)
         );
  OA22X1 U5355 ( .IN1(n6145), .IN2(n5279), .IN3(n5282), .IN4(n6145), .Q(n4425)
         );
  OAI22X1 U5356 ( .IN1(n5342), .IN2(n4426), .IN3(n6454), .IN4(n5343), .QN(
        N10095) );
  OA22X1 U5357 ( .IN1(n5328), .IN2(n4427), .IN3(n6454), .IN4(n5336), .Q(n4426)
         );
  OA22X1 U5358 ( .IN1(n6300), .IN2(n5307), .IN3(n5317), .IN4(n4428), .Q(n4427)
         );
  OA22X1 U5359 ( .IN1(n5293), .IN2(n4429), .IN3(n6300), .IN4(n5301), .Q(n4428)
         );
  OA22X1 U5360 ( .IN1(n6146), .IN2(n5278), .IN3(n5282), .IN4(n6146), .Q(n4429)
         );
  OA22X1 U5362 ( .IN1(n5328), .IN2(n4431), .IN3(n6320), .IN4(n5336), .Q(n4430)
         );
  OA22X1 U5367 ( .IN1(n5328), .IN2(n4435), .IN3(n6321), .IN4(n5336), .Q(n4434)
         );
  OA22X1 U5372 ( .IN1(n5328), .IN2(n4439), .IN3(n6322), .IN4(n5336), .Q(n4438)
         );
  OA22X1 U5377 ( .IN1(n5328), .IN2(n4443), .IN3(n6323), .IN4(n5336), .Q(n4442)
         );
  OA22X1 U5382 ( .IN1(n5328), .IN2(n4447), .IN3(n6324), .IN4(n5336), .Q(n4446)
         );
  OA22X1 U5387 ( .IN1(n5328), .IN2(n4451), .IN3(n6325), .IN4(n5336), .Q(n4450)
         );
  OA22X1 U5392 ( .IN1(n5328), .IN2(n4455), .IN3(n6326), .IN4(n5337), .Q(n4454)
         );
  OA22X1 U5397 ( .IN1(n5328), .IN2(n4459), .IN3(n6327), .IN4(n5337), .Q(n4458)
         );
  OA22X1 U5402 ( .IN1(n5328), .IN2(n4463), .IN3(n6328), .IN4(n5337), .Q(n4462)
         );
  OA22X1 U5407 ( .IN1(n5328), .IN2(n4467), .IN3(n6329), .IN4(n5337), .Q(n4466)
         );
  OA22X1 U5412 ( .IN1(n5328), .IN2(n4471), .IN3(n6330), .IN4(n5337), .Q(n4470)
         );
  OA22X1 U5417 ( .IN1(n5329), .IN2(n4475), .IN3(n6331), .IN4(n5337), .Q(n4474)
         );
  OA22X1 U5422 ( .IN1(n5329), .IN2(n4479), .IN3(n6332), .IN4(n5337), .Q(n4478)
         );
  OA22X1 U5427 ( .IN1(n5329), .IN2(n4483), .IN3(n6333), .IN4(n5337), .Q(n4482)
         );
  OA22X1 U5432 ( .IN1(n5329), .IN2(n4487), .IN3(n6334), .IN4(n5337), .Q(n4486)
         );
  OA22X1 U5437 ( .IN1(n5329), .IN2(n4491), .IN3(n6335), .IN4(n5337), .Q(n4490)
         );
  OA22X1 U5442 ( .IN1(n5329), .IN2(n4495), .IN3(n6336), .IN4(n5337), .Q(n4494)
         );
  OA22X1 U5447 ( .IN1(n5329), .IN2(n4499), .IN3(n6337), .IN4(n5337), .Q(n4498)
         );
  OA22X1 U5452 ( .IN1(n5329), .IN2(n4503), .IN3(n6338), .IN4(n5337), .Q(n4502)
         );
  OA22X1 U5457 ( .IN1(n5329), .IN2(n4507), .IN3(n6339), .IN4(n5337), .Q(n4506)
         );
  OA22X1 U5462 ( .IN1(n5329), .IN2(n4511), .IN3(n6340), .IN4(n5337), .Q(n4510)
         );
  OA22X1 U5467 ( .IN1(n5329), .IN2(n4515), .IN3(n6341), .IN4(n5319), .Q(n4514)
         );
  OA22X1 U5472 ( .IN1(n5329), .IN2(n4519), .IN3(n6342), .IN4(n5320), .Q(n4518)
         );
  OA22X1 U5477 ( .IN1(n5330), .IN2(n4523), .IN3(n6343), .IN4(n5319), .Q(n4522)
         );
  OA22X1 U5482 ( .IN1(n5330), .IN2(n4527), .IN3(n6344), .IN4(n5320), .Q(n4526)
         );
  OA22X1 U5487 ( .IN1(n5330), .IN2(n4531), .IN3(n6345), .IN4(n5319), .Q(n4530)
         );
  OA22X1 U5492 ( .IN1(n5330), .IN2(n4535), .IN3(n6346), .IN4(n5320), .Q(n4534)
         );
  OA22X1 U5497 ( .IN1(n5330), .IN2(n4539), .IN3(n6315), .IN4(n5319), .Q(n4538)
         );
  OA22X1 U5502 ( .IN1(n5330), .IN2(n4543), .IN3(n6316), .IN4(n5320), .Q(n4542)
         );
  OA22X1 U5507 ( .IN1(n5330), .IN2(n4547), .IN3(n6317), .IN4(n5319), .Q(n4546)
         );
  OA22X1 U5512 ( .IN1(n5330), .IN2(n4551), .IN3(n6318), .IN4(n5320), .Q(n4550)
         );
  OA22X1 U5517 ( .IN1(n5330), .IN2(n4555), .IN3(n6319), .IN4(n5319), .Q(n4554)
         );
  OAI22X1 U5521 ( .IN1(n5342), .IN2(n4558), .IN3(n6455), .IN4(n5344), .QN(
        N10062) );
  OA22X1 U5522 ( .IN1(n5330), .IN2(n4559), .IN3(n6455), .IN4(n5320), .Q(n4558)
         );
  OA22X1 U5523 ( .IN1(n6301), .IN2(n5306), .IN3(n5317), .IN4(n4560), .Q(n4559)
         );
  OA22X1 U5524 ( .IN1(n5295), .IN2(n4561), .IN3(n6301), .IN4(n5303), .Q(n4560)
         );
  OA22X1 U5525 ( .IN1(n6147), .IN2(n5278), .IN3(n5282), .IN4(n6147), .Q(n4561)
         );
  OAI22X1 U5526 ( .IN1(n5339), .IN2(n4562), .IN3(n6456), .IN4(n5350), .QN(
        N10061) );
  OA22X1 U5527 ( .IN1(n5330), .IN2(n4563), .IN3(n6456), .IN4(n5319), .Q(n4562)
         );
  OA22X1 U5528 ( .IN1(n6302), .IN2(n5306), .IN3(n5316), .IN4(n4564), .Q(n4563)
         );
  OA22X1 U5529 ( .IN1(n5295), .IN2(n4565), .IN3(n6302), .IN4(n5303), .Q(n4564)
         );
  OA22X1 U5530 ( .IN1(n6148), .IN2(n5278), .IN3(n5282), .IN4(n6148), .Q(n4565)
         );
  OAI22X1 U5531 ( .IN1(n5338), .IN2(n4566), .IN3(n6457), .IN4(n5343), .QN(
        N10060) );
  OA22X1 U5532 ( .IN1(n5330), .IN2(n4567), .IN3(n6457), .IN4(n5320), .Q(n4566)
         );
  OA22X1 U5533 ( .IN1(n6303), .IN2(n5306), .IN3(n5317), .IN4(n4568), .Q(n4567)
         );
  OA22X1 U5534 ( .IN1(n5295), .IN2(n4569), .IN3(n6303), .IN4(n5303), .Q(n4568)
         );
  OA22X1 U5535 ( .IN1(n6149), .IN2(n5278), .IN3(n5282), .IN4(n6149), .Q(n4569)
         );
  OAI22X1 U5536 ( .IN1(n5339), .IN2(n4570), .IN3(n6458), .IN4(n5348), .QN(
        N10059) );
  OA22X1 U5537 ( .IN1(n5322), .IN2(n4571), .IN3(n6458), .IN4(n5320), .Q(n4570)
         );
  OA22X1 U5538 ( .IN1(n6304), .IN2(n5306), .IN3(n5314), .IN4(n4572), .Q(n4571)
         );
  OA22X1 U5539 ( .IN1(n5293), .IN2(n4573), .IN3(n6304), .IN4(n5303), .Q(n4572)
         );
  OA22X1 U5540 ( .IN1(n6150), .IN2(n5278), .IN3(n5282), .IN4(n6150), .Q(n4573)
         );
  OAI22X1 U5541 ( .IN1(n5338), .IN2(n4574), .IN3(n6459), .IN4(n5348), .QN(
        N10058) );
  OA22X1 U5542 ( .IN1(n5321), .IN2(n4575), .IN3(n6459), .IN4(n5320), .Q(n4574)
         );
  OA22X1 U5543 ( .IN1(n6305), .IN2(n5306), .IN3(n5314), .IN4(n4576), .Q(n4575)
         );
  OA22X1 U5544 ( .IN1(n5294), .IN2(n4577), .IN3(n6305), .IN4(n5296), .Q(n4576)
         );
  OA22X1 U5545 ( .IN1(n6151), .IN2(n5278), .IN3(n5282), .IN4(n6151), .Q(n4577)
         );
  NAND4X0 U5546 ( .IN1(n4072), .IN2(n5306), .IN3(n4578), .IN4(n5296), .QN(
        decodedVector_o[3]) );
  NAND4X0 U5547 ( .IN1(n1754), .IN2(decodedPacketValid[4]), .IN3(N2173), .IN4(
        N2172), .QN(n4076) );
  NAND4X0 U5549 ( .IN1(n1752), .IN2(decodedPacketValid[7]), .IN3(N8581), .IN4(
        N8580), .QN(n4070) );
  NAND4X0 U5551 ( .IN1(n1753), .IN2(decodedPacketValid[6]), .IN3(N6445), .IN4(
        N6444), .QN(n4072) );
  OA22X1 U5573 ( .IN1(n5831), .IN2(n4596), .IN3(n5839), .IN4(n5856), .Q(n4595)
         );
  OAI22X1 U5577 ( .IN1(n5846), .IN2(n4599), .IN3(n5852), .IN4(n6384), .QN(
        N10051) );
  OA22X1 U5578 ( .IN1(n5832), .IN2(n4600), .IN3(n5839), .IN4(n6349), .Q(n4599)
         );
  OA22X1 U5579 ( .IN1(n5812), .IN2(n6230), .IN3(n5817), .IN4(n4601), .Q(n4600)
         );
  OA22X1 U5580 ( .IN1(n5796), .IN2(n4602), .IN3(n5801), .IN4(n6195), .Q(n4601)
         );
  OA22X1 U5581 ( .IN1(n5777), .IN2(n6076), .IN3(n5783), .IN4(n6041), .Q(n4602)
         );
  OAI22X1 U5582 ( .IN1(n5846), .IN2(n4603), .IN3(n5852), .IN4(n6376), .QN(
        N10050) );
  OA22X1 U5583 ( .IN1(n5832), .IN2(n4604), .IN3(n5839), .IN4(n6348), .Q(n4603)
         );
  OA22X1 U5584 ( .IN1(n5812), .IN2(n6222), .IN3(n5817), .IN4(n4605), .Q(n4604)
         );
  OA22X1 U5585 ( .IN1(n5796), .IN2(n4606), .IN3(n5802), .IN4(n6194), .Q(n4605)
         );
  OA22X1 U5586 ( .IN1(n5777), .IN2(n6068), .IN3(n5783), .IN4(n6040), .Q(n4606)
         );
  OAI22X1 U5587 ( .IN1(n5846), .IN2(n4607), .IN3(n5852), .IN4(n6373), .QN(
        N10049) );
  OA22X1 U5588 ( .IN1(n5832), .IN2(n4608), .IN3(n5839), .IN4(n6374), .Q(n4607)
         );
  OA22X1 U5589 ( .IN1(n5812), .IN2(n6219), .IN3(n5817), .IN4(n4609), .Q(n4608)
         );
  OA22X1 U5590 ( .IN1(n5796), .IN2(n4610), .IN3(n5802), .IN4(n6220), .Q(n4609)
         );
  OA22X1 U5591 ( .IN1(n5777), .IN2(n6065), .IN3(n5783), .IN4(n6066), .Q(n4610)
         );
  OA22X1 U5593 ( .IN1(n5832), .IN2(n4612), .IN3(n5839), .IN4(n6371), .Q(n4611)
         );
  OAI22X1 U5597 ( .IN1(n5846), .IN2(n4615), .IN3(n5852), .IN4(n6373), .QN(
        N10047) );
  OA22X1 U5598 ( .IN1(n5832), .IN2(n4616), .IN3(n5840), .IN4(n6370), .Q(n4615)
         );
  OA22X1 U5599 ( .IN1(n5812), .IN2(n6219), .IN3(n5817), .IN4(n4617), .Q(n4616)
         );
  OA22X1 U5600 ( .IN1(n5796), .IN2(n4618), .IN3(n5802), .IN4(n6216), .Q(n4617)
         );
  OA22X1 U5601 ( .IN1(n5777), .IN2(n6065), .IN3(n5783), .IN4(n6062), .Q(n4618)
         );
  OAI22X1 U5602 ( .IN1(n5846), .IN2(n4619), .IN3(n5852), .IN4(n6397), .QN(
        N10046) );
  OA22X1 U5603 ( .IN1(n5832), .IN2(n4620), .IN3(n5840), .IN4(n6347), .Q(n4619)
         );
  OA22X1 U5604 ( .IN1(n5812), .IN2(n6245), .IN3(n5817), .IN4(n4621), .Q(n4620)
         );
  OA22X1 U5605 ( .IN1(n5796), .IN2(n4622), .IN3(n5802), .IN4(n6193), .Q(n4621)
         );
  OA22X1 U5606 ( .IN1(n5777), .IN2(n6091), .IN3(n5783), .IN4(n6039), .Q(n4622)
         );
  OAI22X1 U5607 ( .IN1(n5846), .IN2(n4623), .IN3(n5848), .IN4(n5967), .QN(
        N10045) );
  OA22X1 U5608 ( .IN1(n5832), .IN2(n4624), .IN3(n5840), .IN4(n6369), .Q(n4623)
         );
  OA22X1 U5609 ( .IN1(n5812), .IN2(n5952), .IN3(n5818), .IN4(n4625), .Q(n4624)
         );
  OA22X1 U5610 ( .IN1(n5796), .IN2(n4626), .IN3(n5803), .IN4(n6215), .Q(n4625)
         );
  OA22X1 U5611 ( .IN1(n5777), .IN2(n5937), .IN3(n5784), .IN4(n6061), .Q(n4626)
         );
  OAI22X1 U5612 ( .IN1(n5846), .IN2(n4627), .IN3(n5851), .IN4(n5968), .QN(
        N10044) );
  OA22X1 U5613 ( .IN1(n5832), .IN2(n4628), .IN3(n5840), .IN4(n6368), .Q(n4627)
         );
  OA22X1 U5614 ( .IN1(n5812), .IN2(n5953), .IN3(n5818), .IN4(n4629), .Q(n4628)
         );
  OA22X1 U5615 ( .IN1(n5796), .IN2(n4630), .IN3(n5803), .IN4(n6214), .Q(n4629)
         );
  OA22X1 U5616 ( .IN1(n5777), .IN2(n5938), .IN3(n5784), .IN4(n6060), .Q(n4630)
         );
  OAI22X1 U5617 ( .IN1(n5846), .IN2(n4631), .IN3(n5852), .IN4(n5969), .QN(
        N10043) );
  OA22X1 U5618 ( .IN1(n5832), .IN2(n4632), .IN3(n5840), .IN4(n6367), .Q(n4631)
         );
  OA22X1 U5619 ( .IN1(n5812), .IN2(n5954), .IN3(n5818), .IN4(n4633), .Q(n4632)
         );
  OA22X1 U5620 ( .IN1(n5796), .IN2(n4634), .IN3(n5803), .IN4(n6213), .Q(n4633)
         );
  OA22X1 U5621 ( .IN1(n5777), .IN2(n5939), .IN3(n5784), .IN4(n6059), .Q(n4634)
         );
  OAI22X1 U5622 ( .IN1(n5847), .IN2(n4635), .IN3(n5850), .IN4(n5970), .QN(
        N10042) );
  OA22X1 U5623 ( .IN1(n5832), .IN2(n4636), .IN3(n5841), .IN4(n6366), .Q(n4635)
         );
  OA22X1 U5624 ( .IN1(n5812), .IN2(n5955), .IN3(n5818), .IN4(n4637), .Q(n4636)
         );
  OA22X1 U5625 ( .IN1(n5796), .IN2(n4638), .IN3(n5803), .IN4(n6212), .Q(n4637)
         );
  OA22X1 U5626 ( .IN1(n5777), .IN2(n5940), .IN3(n5784), .IN4(n6058), .Q(n4638)
         );
  OAI22X1 U5627 ( .IN1(n5847), .IN2(n4639), .IN3(n5853), .IN4(n5971), .QN(
        N10041) );
  OA22X1 U5628 ( .IN1(n5832), .IN2(n4640), .IN3(n5841), .IN4(n6365), .Q(n4639)
         );
  OA22X1 U5629 ( .IN1(n5812), .IN2(n5956), .IN3(n5818), .IN4(n4641), .Q(n4640)
         );
  OA22X1 U5630 ( .IN1(n5796), .IN2(n4642), .IN3(n5803), .IN4(n6211), .Q(n4641)
         );
  OA22X1 U5631 ( .IN1(n5777), .IN2(n5941), .IN3(n5784), .IN4(n6057), .Q(n4642)
         );
  OAI22X1 U5632 ( .IN1(n5847), .IN2(n4643), .IN3(n5853), .IN4(n5972), .QN(
        N10040) );
  OA22X1 U5633 ( .IN1(n5832), .IN2(n4644), .IN3(n5841), .IN4(n6364), .Q(n4643)
         );
  OA22X1 U5634 ( .IN1(n5812), .IN2(n5957), .IN3(n5816), .IN4(n4645), .Q(n4644)
         );
  OA22X1 U5635 ( .IN1(n5796), .IN2(n4646), .IN3(n5804), .IN4(n6210), .Q(n4645)
         );
  OA22X1 U5636 ( .IN1(n5777), .IN2(n5942), .IN3(n5784), .IN4(n6056), .Q(n4646)
         );
  OAI22X1 U5637 ( .IN1(n5847), .IN2(n4647), .IN3(n5853), .IN4(n5973), .QN(
        N10039) );
  OA22X1 U5638 ( .IN1(n5833), .IN2(n4648), .IN3(n5841), .IN4(n6363), .Q(n4647)
         );
  OA22X1 U5639 ( .IN1(n5812), .IN2(n5958), .IN3(n5817), .IN4(n4649), .Q(n4648)
         );
  OA22X1 U5640 ( .IN1(n5797), .IN2(n4650), .IN3(n5804), .IN4(n6209), .Q(n4649)
         );
  OA22X1 U5641 ( .IN1(n5777), .IN2(n5943), .IN3(n5782), .IN4(n6055), .Q(n4650)
         );
  OAI22X1 U5642 ( .IN1(n5847), .IN2(n4651), .IN3(n5853), .IN4(n5974), .QN(
        N10038) );
  OA22X1 U5643 ( .IN1(n5833), .IN2(n4652), .IN3(n5841), .IN4(n6362), .Q(n4651)
         );
  OA22X1 U5644 ( .IN1(n5812), .IN2(n5959), .IN3(n5821), .IN4(n4653), .Q(n4652)
         );
  OA22X1 U5645 ( .IN1(n5797), .IN2(n4654), .IN3(n5804), .IN4(n6208), .Q(n4653)
         );
  OA22X1 U5646 ( .IN1(n5777), .IN2(n5944), .IN3(n5786), .IN4(n6054), .Q(n4654)
         );
  OAI22X1 U5647 ( .IN1(n5847), .IN2(n4655), .IN3(n5853), .IN4(n5975), .QN(
        N10037) );
  OA22X1 U5648 ( .IN1(n5833), .IN2(n4656), .IN3(n5842), .IN4(n6308), .Q(n4655)
         );
  OA22X1 U5649 ( .IN1(n5812), .IN2(n5960), .IN3(n5820), .IN4(n4657), .Q(n4656)
         );
  OA22X1 U5650 ( .IN1(n5797), .IN2(n4658), .IN3(n5804), .IN4(n6154), .Q(n4657)
         );
  OA22X1 U5651 ( .IN1(n5777), .IN2(n5945), .IN3(n5782), .IN4(n6000), .Q(n4658)
         );
  OAI22X1 U5652 ( .IN1(n5847), .IN2(n4659), .IN3(n5848), .IN4(n5976), .QN(
        N10036) );
  OA22X1 U5653 ( .IN1(n5833), .IN2(n4660), .IN3(n5842), .IN4(n6309), .Q(n4659)
         );
  OA22X1 U5654 ( .IN1(n5812), .IN2(n5961), .IN3(n5818), .IN4(n4661), .Q(n4660)
         );
  OA22X1 U5655 ( .IN1(n5797), .IN2(n4662), .IN3(n5804), .IN4(n6155), .Q(n4661)
         );
  OA22X1 U5656 ( .IN1(n5777), .IN2(n5946), .IN3(n5781), .IN4(n6001), .Q(n4662)
         );
  OAI22X1 U5657 ( .IN1(n5847), .IN2(n4663), .IN3(n5852), .IN4(n5977), .QN(
        N10035) );
  OA22X1 U5658 ( .IN1(n5833), .IN2(n4664), .IN3(n5842), .IN4(n6310), .Q(n4663)
         );
  OA22X1 U5659 ( .IN1(n5812), .IN2(n5962), .IN3(n5815), .IN4(n4665), .Q(n4664)
         );
  OA22X1 U5660 ( .IN1(n5797), .IN2(n4666), .IN3(n5805), .IN4(n6156), .Q(n4665)
         );
  OA22X1 U5661 ( .IN1(n5777), .IN2(n5947), .IN3(n5780), .IN4(n6002), .Q(n4666)
         );
  OAI22X1 U5662 ( .IN1(n5847), .IN2(n4667), .IN3(n5853), .IN4(n5978), .QN(
        N10034) );
  OA22X1 U5663 ( .IN1(n5833), .IN2(n4668), .IN3(n5842), .IN4(n6311), .Q(n4667)
         );
  OA22X1 U5664 ( .IN1(n5812), .IN2(n5963), .IN3(n5820), .IN4(n4669), .Q(n4668)
         );
  OA22X1 U5665 ( .IN1(n5797), .IN2(n4670), .IN3(n5805), .IN4(n6157), .Q(n4669)
         );
  OA22X1 U5666 ( .IN1(n5777), .IN2(n5948), .IN3(n5782), .IN4(n6003), .Q(n4670)
         );
  OAI22X1 U5667 ( .IN1(n5847), .IN2(n4671), .IN3(n5853), .IN4(n5979), .QN(
        N10033) );
  OA22X1 U5668 ( .IN1(n5833), .IN2(n4672), .IN3(n5842), .IN4(n6312), .Q(n4671)
         );
  OA22X1 U5669 ( .IN1(n5812), .IN2(n5964), .IN3(n5814), .IN4(n4673), .Q(n4672)
         );
  OA22X1 U5670 ( .IN1(n5797), .IN2(n4674), .IN3(n5805), .IN4(n6158), .Q(n4673)
         );
  OA22X1 U5671 ( .IN1(n5777), .IN2(n5949), .IN3(n5783), .IN4(n6004), .Q(n4674)
         );
  OAI22X1 U5672 ( .IN1(n5847), .IN2(n4675), .IN3(n5848), .IN4(n5980), .QN(
        N10032) );
  OA22X1 U5673 ( .IN1(n5833), .IN2(n4676), .IN3(n5840), .IN4(n6313), .Q(n4675)
         );
  OA22X1 U5674 ( .IN1(n5812), .IN2(n5965), .IN3(n5815), .IN4(n4677), .Q(n4676)
         );
  OA22X1 U5675 ( .IN1(n5797), .IN2(n4678), .IN3(n5805), .IN4(n6159), .Q(n4677)
         );
  OA22X1 U5676 ( .IN1(n5777), .IN2(n5950), .IN3(n5780), .IN4(n6005), .Q(n4678)
         );
  OAI22X1 U5677 ( .IN1(n5847), .IN2(n4679), .IN3(n5852), .IN4(n5981), .QN(
        N10031) );
  OA22X1 U5678 ( .IN1(n5833), .IN2(n4680), .IN3(n5841), .IN4(n6314), .Q(n4679)
         );
  OA22X1 U5679 ( .IN1(n5812), .IN2(n5966), .IN3(n5818), .IN4(n4681), .Q(n4680)
         );
  OA22X1 U5680 ( .IN1(n5797), .IN2(n4682), .IN3(n5805), .IN4(n6160), .Q(n4681)
         );
  OA22X1 U5681 ( .IN1(n5777), .IN2(n5951), .IN3(n5779), .IN4(n6006), .Q(n4682)
         );
  OAI22X1 U5682 ( .IN1(n5847), .IN2(n4683), .IN3(n5849), .IN4(n6375), .QN(
        N10030) );
  OA22X1 U5683 ( .IN1(n5833), .IN2(n4684), .IN3(n5842), .IN4(n6307), .Q(n4683)
         );
  OA22X1 U5684 ( .IN1(n5812), .IN2(n6221), .IN3(n5819), .IN4(n4685), .Q(n4684)
         );
  OA22X1 U5685 ( .IN1(n5797), .IN2(n4686), .IN3(n5805), .IN4(n6153), .Q(n4685)
         );
  OA22X1 U5686 ( .IN1(n5777), .IN2(n6067), .IN3(n5781), .IN4(n5999), .Q(n4686)
         );
  OAI22X1 U5687 ( .IN1(n5847), .IN2(n4687), .IN3(n5853), .IN4(n6372), .QN(
        N10028) );
  OA22X1 U5688 ( .IN1(n5833), .IN2(n4688), .IN3(n5836), .IN4(n6306), .Q(n4687)
         );
  OA22X1 U5689 ( .IN1(n5812), .IN2(n6218), .IN3(n5819), .IN4(n4689), .Q(n4688)
         );
  OA22X1 U5690 ( .IN1(n5797), .IN2(n4690), .IN3(n5789), .IN4(n6152), .Q(n4689)
         );
  OA22X1 U5691 ( .IN1(n5777), .IN2(n6064), .IN3(n5780), .IN4(n5998), .Q(n4690)
         );
  NAND4X0 U5692 ( .IN1(n828), .IN2(n5810), .IN3(n4691), .IN4(n4692), .QN(
        decodedVector_o[2]) );
  AND3X1 U5693 ( .IN1(n5778), .IN2(n826), .IN3(n832), .Q(n4692) );
  OAI22X1 U5694 ( .IN1(n5847), .IN2(n4693), .IN3(n5849), .IN4(n6377), .QN(
        N10026) );
  OA22X1 U5695 ( .IN1(n5833), .IN2(n4694), .IN3(n5825), .IN4(n6422), .Q(n4693)
         );
  OA22X1 U5696 ( .IN1(n5812), .IN2(n6223), .IN3(n5819), .IN4(n4695), .Q(n4694)
         );
  OA22X1 U5697 ( .IN1(n5797), .IN2(n4696), .IN3(n5788), .IN4(n6268), .Q(n4695)
         );
  OA22X1 U5698 ( .IN1(n5777), .IN2(n6069), .IN3(n5779), .IN4(n6114), .Q(n4696)
         );
  OAI22X1 U5699 ( .IN1(n5847), .IN2(n4697), .IN3(n826), .IN4(n6378), .QN(
        N10025) );
  OA22X1 U5700 ( .IN1(n5834), .IN2(n4698), .IN3(n5839), .IN4(n6421), .Q(n4697)
         );
  OA22X1 U5701 ( .IN1(n5812), .IN2(n6224), .IN3(n5819), .IN4(n4699), .Q(n4698)
         );
  OA22X1 U5702 ( .IN1(n5798), .IN2(n4700), .IN3(n5787), .IN4(n6267), .Q(n4699)
         );
  OA22X1 U5703 ( .IN1(n5777), .IN2(n6070), .IN3(n5785), .IN4(n6113), .Q(n4700)
         );
  OAI22X1 U5704 ( .IN1(n5847), .IN2(n4701), .IN3(n5853), .IN4(n6379), .QN(
        N10024) );
  OA22X1 U5705 ( .IN1(n5834), .IN2(n4702), .IN3(n5824), .IN4(n6420), .Q(n4701)
         );
  OA22X1 U5706 ( .IN1(n5812), .IN2(n6225), .IN3(n5819), .IN4(n4703), .Q(n4702)
         );
  OA22X1 U5707 ( .IN1(n5798), .IN2(n4704), .IN3(n5806), .IN4(n6266), .Q(n4703)
         );
  OA22X1 U5708 ( .IN1(n5777), .IN2(n6071), .IN3(n5784), .IN4(n6112), .Q(n4704)
         );
  OAI22X1 U5709 ( .IN1(n5847), .IN2(n4705), .IN3(n826), .IN4(n6380), .QN(
        N10023) );
  OA22X1 U5710 ( .IN1(n5834), .IN2(n4706), .IN3(n5825), .IN4(n6419), .Q(n4705)
         );
  OA22X1 U5711 ( .IN1(n5812), .IN2(n6226), .IN3(n5820), .IN4(n4707), .Q(n4706)
         );
  OA22X1 U5712 ( .IN1(n5798), .IN2(n4708), .IN3(n5806), .IN4(n6265), .Q(n4707)
         );
  OA22X1 U5713 ( .IN1(n5777), .IN2(n6072), .IN3(n5785), .IN4(n6111), .Q(n4708)
         );
  OAI22X1 U5714 ( .IN1(n5847), .IN2(n4709), .IN3(n5851), .IN4(n6381), .QN(
        N10022) );
  OA22X1 U5715 ( .IN1(n5834), .IN2(n4710), .IN3(n5839), .IN4(n6418), .Q(n4709)
         );
  OA22X1 U5716 ( .IN1(n5812), .IN2(n6227), .IN3(n5818), .IN4(n4711), .Q(n4710)
         );
  OA22X1 U5717 ( .IN1(n5798), .IN2(n4712), .IN3(n5806), .IN4(n6264), .Q(n4711)
         );
  OA22X1 U5718 ( .IN1(n5777), .IN2(n6073), .IN3(n5784), .IN4(n6110), .Q(n4712)
         );
  OAI22X1 U5719 ( .IN1(n5847), .IN2(n4713), .IN3(n5850), .IN4(n6382), .QN(
        N10021) );
  OA22X1 U5720 ( .IN1(n5834), .IN2(n4714), .IN3(n5822), .IN4(n6417), .Q(n4713)
         );
  OA22X1 U5721 ( .IN1(n5813), .IN2(n6228), .IN3(n5821), .IN4(n4715), .Q(n4714)
         );
  OA22X1 U5722 ( .IN1(n5798), .IN2(n4716), .IN3(n5806), .IN4(n6263), .Q(n4715)
         );
  OA22X1 U5723 ( .IN1(n5777), .IN2(n6074), .IN3(n5786), .IN4(n6109), .Q(n4716)
         );
  OAI22X1 U5724 ( .IN1(n5847), .IN2(n4717), .IN3(n5850), .IN4(n6383), .QN(
        N10020) );
  OA22X1 U5725 ( .IN1(n5834), .IN2(n4718), .IN3(n5825), .IN4(n6416), .Q(n4717)
         );
  OA22X1 U5726 ( .IN1(n5813), .IN2(n6229), .IN3(n5821), .IN4(n4719), .Q(n4718)
         );
  OA22X1 U5727 ( .IN1(n5798), .IN2(n4720), .IN3(n5806), .IN4(n6262), .Q(n4719)
         );
  OA22X1 U5728 ( .IN1(n5778), .IN2(n6075), .IN3(n5783), .IN4(n6108), .Q(n4720)
         );
  OAI22X1 U5729 ( .IN1(n5847), .IN2(n4721), .IN3(n5850), .IN4(n6385), .QN(
        N10019) );
  OA22X1 U5730 ( .IN1(n5834), .IN2(n4722), .IN3(n5822), .IN4(n6359), .Q(n4721)
         );
  OA22X1 U5731 ( .IN1(n5813), .IN2(n6231), .IN3(n5819), .IN4(n4723), .Q(n4722)
         );
  OA22X1 U5732 ( .IN1(n5798), .IN2(n4724), .IN3(n5806), .IN4(n6205), .Q(n4723)
         );
  OA22X1 U5733 ( .IN1(n5778), .IN2(n6077), .IN3(n5783), .IN4(n6051), .Q(n4724)
         );
  OAI22X1 U5734 ( .IN1(n5847), .IN2(n4725), .IN3(n5848), .IN4(n6386), .QN(
        N10018) );
  OA22X1 U5735 ( .IN1(n5834), .IN2(n4726), .IN3(n5823), .IN4(n6358), .Q(n4725)
         );
  OA22X1 U5736 ( .IN1(n5813), .IN2(n6232), .IN3(n5820), .IN4(n4727), .Q(n4726)
         );
  OA22X1 U5737 ( .IN1(n5798), .IN2(n4728), .IN3(n5807), .IN4(n6204), .Q(n4727)
         );
  OA22X1 U5738 ( .IN1(n5778), .IN2(n6078), .IN3(n5785), .IN4(n6050), .Q(n4728)
         );
  OAI22X1 U5739 ( .IN1(n5847), .IN2(n4729), .IN3(n5853), .IN4(n6387), .QN(
        N10017) );
  OA22X1 U5740 ( .IN1(n5834), .IN2(n4730), .IN3(n5824), .IN4(n6357), .Q(n4729)
         );
  OA22X1 U5741 ( .IN1(n5813), .IN2(n6233), .IN3(n5820), .IN4(n4731), .Q(n4730)
         );
  OA22X1 U5742 ( .IN1(n5798), .IN2(n4732), .IN3(n5807), .IN4(n6203), .Q(n4731)
         );
  OA22X1 U5743 ( .IN1(n5778), .IN2(n6079), .IN3(n5785), .IN4(n6049), .Q(n4732)
         );
  OAI22X1 U5744 ( .IN1(n5847), .IN2(n4733), .IN3(n5850), .IN4(n6388), .QN(
        N10016) );
  OA22X1 U5745 ( .IN1(n5834), .IN2(n4734), .IN3(n5837), .IN4(n6356), .Q(n4733)
         );
  OA22X1 U5746 ( .IN1(n5813), .IN2(n6234), .IN3(n5820), .IN4(n4735), .Q(n4734)
         );
  OA22X1 U5747 ( .IN1(n5798), .IN2(n4736), .IN3(n5807), .IN4(n6202), .Q(n4735)
         );
  OA22X1 U5748 ( .IN1(n5778), .IN2(n6080), .IN3(n5785), .IN4(n6048), .Q(n4736)
         );
  OAI22X1 U5749 ( .IN1(n5847), .IN2(n4737), .IN3(n5849), .IN4(n6389), .QN(
        N10015) );
  OA22X1 U5750 ( .IN1(n5834), .IN2(n4738), .IN3(n5842), .IN4(n6355), .Q(n4737)
         );
  OA22X1 U5751 ( .IN1(n5813), .IN2(n6235), .IN3(n5820), .IN4(n4739), .Q(n4738)
         );
  OA22X1 U5752 ( .IN1(n5798), .IN2(n4740), .IN3(n5807), .IN4(n6201), .Q(n4739)
         );
  OA22X1 U5753 ( .IN1(n5778), .IN2(n6081), .IN3(n5785), .IN4(n6047), .Q(n4740)
         );
  OAI22X1 U5754 ( .IN1(n5847), .IN2(n4741), .IN3(n5853), .IN4(n6390), .QN(
        N10014) );
  OA22X1 U5755 ( .IN1(n5834), .IN2(n4742), .IN3(n5838), .IN4(n6354), .Q(n4741)
         );
  OA22X1 U5756 ( .IN1(n5813), .IN2(n6236), .IN3(n5820), .IN4(n4743), .Q(n4742)
         );
  OA22X1 U5757 ( .IN1(n5798), .IN2(n4744), .IN3(n5800), .IN4(n6200), .Q(n4743)
         );
  OA22X1 U5758 ( .IN1(n5778), .IN2(n6082), .IN3(n5785), .IN4(n6046), .Q(n4744)
         );
  OAI22X1 U5759 ( .IN1(n5847), .IN2(n4745), .IN3(n5849), .IN4(n6391), .QN(
        N10013) );
  OA22X1 U5760 ( .IN1(n5835), .IN2(n4746), .IN3(n5841), .IN4(n6353), .Q(n4745)
         );
  OA22X1 U5761 ( .IN1(n5813), .IN2(n6237), .IN3(n5821), .IN4(n4747), .Q(n4746)
         );
  OA22X1 U5762 ( .IN1(n5799), .IN2(n4748), .IN3(n5807), .IN4(n6199), .Q(n4747)
         );
  OA22X1 U5763 ( .IN1(n5778), .IN2(n6083), .IN3(n5786), .IN4(n6045), .Q(n4748)
         );
  OAI22X1 U5764 ( .IN1(n5847), .IN2(n4749), .IN3(n5853), .IN4(n6400), .QN(
        N10012) );
  OA22X1 U5765 ( .IN1(n5835), .IN2(n4750), .IN3(n5836), .IN4(n6415), .Q(n4749)
         );
  OA22X1 U5766 ( .IN1(n5813), .IN2(n6246), .IN3(n5821), .IN4(n4751), .Q(n4750)
         );
  OA22X1 U5767 ( .IN1(n5799), .IN2(n4752), .IN3(n5801), .IN4(n6261), .Q(n4751)
         );
  OA22X1 U5768 ( .IN1(n5778), .IN2(n6092), .IN3(n5786), .IN4(n6107), .Q(n4752)
         );
  OAI22X1 U5769 ( .IN1(n5847), .IN2(n4753), .IN3(n5851), .IN4(n6406), .QN(
        N10011) );
  OA22X1 U5770 ( .IN1(n5835), .IN2(n4754), .IN3(n5822), .IN4(n6414), .Q(n4753)
         );
  OA22X1 U5771 ( .IN1(n5813), .IN2(n6252), .IN3(n5821), .IN4(n4755), .Q(n4754)
         );
  OA22X1 U5772 ( .IN1(n5799), .IN2(n4756), .IN3(n5801), .IN4(n6260), .Q(n4755)
         );
  OA22X1 U5773 ( .IN1(n5778), .IN2(n6098), .IN3(n5786), .IN4(n6106), .Q(n4756)
         );
  OAI22X1 U5774 ( .IN1(n5847), .IN2(n4757), .IN3(n826), .IN4(n6407), .QN(
        N10010) );
  OA22X1 U5775 ( .IN1(n5835), .IN2(n4758), .IN3(n5823), .IN4(n6413), .Q(n4757)
         );
  OA22X1 U5776 ( .IN1(n5813), .IN2(n6253), .IN3(n5821), .IN4(n4759), .Q(n4758)
         );
  OA22X1 U5777 ( .IN1(n5799), .IN2(n4760), .IN3(n5802), .IN4(n6259), .Q(n4759)
         );
  OA22X1 U5778 ( .IN1(n5778), .IN2(n6099), .IN3(n5786), .IN4(n6105), .Q(n4760)
         );
  OAI22X1 U5779 ( .IN1(n5847), .IN2(n4761), .IN3(n5848), .IN4(n6408), .QN(
        N10009) );
  OA22X1 U5780 ( .IN1(n5835), .IN2(n4762), .IN3(n5824), .IN4(n6412), .Q(n4761)
         );
  OA22X1 U5781 ( .IN1(n5813), .IN2(n6254), .IN3(n5821), .IN4(n4763), .Q(n4762)
         );
  OA22X1 U5782 ( .IN1(n5799), .IN2(n4764), .IN3(n5789), .IN4(n6258), .Q(n4763)
         );
  OA22X1 U5783 ( .IN1(n5778), .IN2(n6100), .IN3(n5786), .IN4(n6104), .Q(n4764)
         );
  OAI22X1 U5784 ( .IN1(n5847), .IN2(n4765), .IN3(n826), .IN4(n6409), .QN(
        N10008) );
  OA22X1 U5785 ( .IN1(n5835), .IN2(n4766), .IN3(n5837), .IN4(n6411), .Q(n4765)
         );
  OA22X1 U5786 ( .IN1(n5813), .IN2(n6255), .IN3(n5816), .IN4(n4767), .Q(n4766)
         );
  OA22X1 U5787 ( .IN1(n5799), .IN2(n4768), .IN3(n5788), .IN4(n6257), .Q(n4767)
         );
  OA22X1 U5788 ( .IN1(n5778), .IN2(n6101), .IN3(n5782), .IN4(n6103), .Q(n4768)
         );
  OAI22X1 U5789 ( .IN1(n5847), .IN2(n4769), .IN3(n5851), .IN4(n6401), .QN(
        N10007) );
  OA22X1 U5790 ( .IN1(n5835), .IN2(n4770), .IN3(n5838), .IN4(n6410), .Q(n4769)
         );
  OA22X1 U5791 ( .IN1(n5813), .IN2(n6247), .IN3(n5818), .IN4(n4771), .Q(n4770)
         );
  OA22X1 U5792 ( .IN1(n5799), .IN2(n4772), .IN3(n5804), .IN4(n6256), .Q(n4771)
         );
  OA22X1 U5793 ( .IN1(n5778), .IN2(n6093), .IN3(n5785), .IN4(n6102), .Q(n4772)
         );
  OAI22X1 U5794 ( .IN1(n5847), .IN2(n4773), .IN3(n5850), .IN4(n6399), .QN(
        N10006) );
  OA22X1 U5795 ( .IN1(n5835), .IN2(n4774), .IN3(n5840), .IN4(n6352), .Q(n4773)
         );
  OA22X1 U5796 ( .IN1(n5813), .IN2(n6244), .IN3(n5821), .IN4(n4775), .Q(n4774)
         );
  OA22X1 U5797 ( .IN1(n5799), .IN2(n4776), .IN3(n5801), .IN4(n6198), .Q(n4775)
         );
  OA22X1 U5798 ( .IN1(n5778), .IN2(n6090), .IN3(n5784), .IN4(n6044), .Q(n4776)
         );
  OAI22X1 U5799 ( .IN1(n5847), .IN2(n4777), .IN3(n5848), .IN4(n6398), .QN(
        N10005) );
  OA22X1 U5800 ( .IN1(n5835), .IN2(n4778), .IN3(n5822), .IN4(n6402), .Q(n4777)
         );
  OA22X1 U5801 ( .IN1(n5813), .IN2(n6243), .IN3(n5817), .IN4(n4779), .Q(n4778)
         );
  OA22X1 U5802 ( .IN1(n5799), .IN2(n4780), .IN3(n5803), .IN4(n6248), .Q(n4779)
         );
  OA22X1 U5803 ( .IN1(n5778), .IN2(n6089), .IN3(n5786), .IN4(n6094), .Q(n4780)
         );
  OAI22X1 U5804 ( .IN1(n5847), .IN2(n4781), .IN3(n5849), .IN4(n6397), .QN(
        N10004) );
  OA22X1 U5805 ( .IN1(n5835), .IN2(n4782), .IN3(n5824), .IN4(n6403), .Q(n4781)
         );
  OA22X1 U5806 ( .IN1(n5813), .IN2(n6242), .IN3(n5816), .IN4(n4783), .Q(n4782)
         );
  OA22X1 U5807 ( .IN1(n5799), .IN2(n4784), .IN3(n5805), .IN4(n6249), .Q(n4783)
         );
  OA22X1 U5808 ( .IN1(n5778), .IN2(n6090), .IN3(n5785), .IN4(n6095), .Q(n4784)
         );
  OAI22X1 U5809 ( .IN1(n5847), .IN2(n4785), .IN3(n5850), .IN4(n6396), .QN(
        N10003) );
  OA22X1 U5810 ( .IN1(n5835), .IN2(n4786), .IN3(n5823), .IN4(n6404), .Q(n4785)
         );
  OA22X1 U5811 ( .IN1(n5813), .IN2(n6241), .IN3(n5819), .IN4(n4787), .Q(n4786)
         );
  OA22X1 U5812 ( .IN1(n5799), .IN2(n4788), .IN3(n5802), .IN4(n6250), .Q(n4787)
         );
  OA22X1 U5813 ( .IN1(n5778), .IN2(n6088), .IN3(n5780), .IN4(n6096), .Q(n4788)
         );
  OAI22X1 U5814 ( .IN1(n5847), .IN2(n4789), .IN3(n826), .IN4(n6395), .QN(
        N10002) );
  OA22X1 U5815 ( .IN1(n5835), .IN2(n4790), .IN3(n5837), .IN4(n6405), .Q(n4789)
         );
  OA22X1 U5816 ( .IN1(n5813), .IN2(n6244), .IN3(n5819), .IN4(n4791), .Q(n4790)
         );
  OA22X1 U5817 ( .IN1(n5799), .IN2(n4792), .IN3(n5806), .IN4(n6251), .Q(n4791)
         );
  OA22X1 U5818 ( .IN1(n5778), .IN2(n6087), .IN3(n5786), .IN4(n6097), .Q(n4792)
         );
  OAI22X1 U5819 ( .IN1(n5847), .IN2(n4793), .IN3(n5851), .IN4(n6394), .QN(
        N10001) );
  OA22X1 U5820 ( .IN1(n5829), .IN2(n4794), .IN3(n5838), .IN4(n6393), .Q(n4793)
         );
  OA22X1 U5821 ( .IN1(n5813), .IN2(n6240), .IN3(n5816), .IN4(n4795), .Q(n4794)
         );
  OA22X1 U5822 ( .IN1(n5794), .IN2(n4796), .IN3(n5807), .IN4(n6239), .Q(n4795)
         );
  OA22X1 U5823 ( .IN1(n5778), .IN2(n6086), .IN3(n5782), .IN4(n6085), .Q(n4796)
         );
  OAI22X1 U5824 ( .IN1(n5843), .IN2(n4797), .IN3(n826), .IN4(n6361), .QN(
        N10000) );
  OA22X1 U5825 ( .IN1(n5830), .IN2(n4798), .IN3(n5840), .IN4(n6360), .Q(n4797)
         );
  OA22X1 U5826 ( .IN1(n5810), .IN2(n6207), .IN3(n5821), .IN4(n4799), .Q(n4798)
         );
  OA22X1 U5827 ( .IN1(n5793), .IN2(n4800), .IN3(n5801), .IN4(n6206), .Q(n4799)
         );
  OA22X1 U5828 ( .IN1(n5775), .IN2(n6053), .IN3(n5782), .IN4(n6052), .Q(n4800)
         );
  NAND4X0 U5835 ( .IN1(n1754), .IN2(decodedPacketValid[4]), .IN3(N2173), .IN4(
        n5995), .QN(n832) );
  NAND4X0 U5847 ( .IN1(n1753), .IN2(decodedPacketValid[6]), .IN3(N6445), .IN4(
        n5993), .QN(n828) );
  NAND4X0 U5853 ( .IN1(n1752), .IN2(decodedPacketValid[7]), .IN3(N8581), .IN4(
        n5992), .QN(n826) );
  NOR3X0 U5858 ( .IN1(N8583), .IN2(N8585), .IN3(N8584), .QN(n4837) );
  Decode_PISA_0 decode0_PISA ( .instPacketValid_i(inst0PacketValid_i), 
        .instPacket_i(inst0Packet_i), .decodedPacket0Valid_o(N389), 
        .decodedPacket0_o({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        \decodedPacket[0][121] , \decodedPacket[0][120] , 
        \decodedPacket[0][119] , \decodedPacket[0][118] , 
        \decodedPacket[0][117] , \decodedPacket[0][116] , 
        \decodedPacket[0][115] , \decodedPacket[0][114] , 
        \decodedPacket[0][113] , \decodedPacket[0][112] , 
        \decodedPacket[0][111] , \decodedPacket[0][110] , 
        \decodedPacket[0][109] , \decodedPacket[0][108] , 
        \decodedPacket[0][107] , \decodedPacket[0][106] , 
        \decodedPacket[0][105] , \decodedPacket[0][104] , 
        \decodedPacket[0][103] , \decodedPacket[0][102] , 
        \decodedPacket[0][101] , \decodedPacket[0][100] , 
        \decodedPacket[0][99] , \decodedPacket[0][98] , \decodedPacket[0][97] , 
        \decodedPacket[0][96] , \decodedPacket[0][95] , \decodedPacket[0][94] , 
        \decodedPacket[0][93] , \decodedPacket[0][92] , \decodedPacket[0][91] , 
        \decodedPacket[0][90] , \decodedPacket[0][89] , \decodedPacket[0][88] , 
        \decodedPacket[0][87] , \decodedPacket[0][86] , \decodedPacket[0][85] , 
        \decodedPacket[0][84] , \decodedPacket[0][83] , \decodedPacket[0][82] , 
        \decodedPacket[0][81] , \decodedPacket[0][80] , \decodedPacket[0][79] , 
        \decodedPacket[0][78] , \decodedPacket[0][77] , \decodedPacket[0][76] , 
        \decodedPacket[0][75] , \decodedPacket[0][74] , \decodedPacket[0][73] , 
        \decodedPacket[0][72] , \decodedPacket[0][71] , \decodedPacket[0][70] , 
        \decodedPacket[0][69] , \decodedPacket[0][68] , \decodedPacket[0][67] , 
        \decodedPacket[0][66] , \decodedPacket[0][65] , \decodedPacket[0][64] , 
        \decodedPacket[0][63] , \decodedPacket[0][62] , \decodedPacket[0][61] , 
        \decodedPacket[0][60] , \decodedPacket[0][59] , \decodedPacket[0][58] , 
        \decodedPacket[0][57] , \decodedPacket[0][56] , \decodedPacket[0][55] , 
        \decodedPacket[0][54] , \decodedPacket[0][53] , \decodedPacket[0][52] , 
        \decodedPacket[0][51] , \decodedPacket[0][50] , \decodedPacket[0][49] , 
        \decodedPacket[0][48] , \decodedPacket[0][47] , \decodedPacket[0][46] , 
        \decodedPacket[0][45] , \decodedPacket[0][44] , \decodedPacket[0][43] , 
        \decodedPacket[0][42] , \decodedPacket[0][41] , \decodedPacket[0][40] , 
        \decodedPacket[0][39] , \decodedPacket[0][38] , \decodedPacket[0][37] , 
        \decodedPacket[0][36] , \decodedPacket[0][35] , \decodedPacket[0][34] , 
        \decodedPacket[0][33] , \decodedPacket[0][32] , \decodedPacket[0][31] , 
        \decodedPacket[0][30] , \decodedPacket[0][29] , \decodedPacket[0][28] , 
        \decodedPacket[0][27] , \decodedPacket[0][26] , \decodedPacket[0][25] , 
        \decodedPacket[0][24] , \decodedPacket[0][23] , \decodedPacket[0][22] , 
        \decodedPacket[0][21] , \decodedPacket[0][20] , \decodedPacket[0][19] , 
        \decodedPacket[0][18] , \decodedPacket[0][17] , \decodedPacket[0][16] , 
        \decodedPacket[0][15] , \decodedPacket[0][14] , \decodedPacket[0][13] , 
        \decodedPacket[0][12] , \decodedPacket[0][11] , \decodedPacket[0][10] , 
        \decodedPacket[0][9] , \decodedPacket[0][8] , \decodedPacket[0][7] , 
        \decodedPacket[0][6] , \decodedPacket[0][5] , \decodedPacket[0][4] , 
        \decodedPacket[0][3] , \decodedPacket[0][2] , \decodedPacket[0][1] , 
        \decodedPacket[0][0] }), .decodedPacket1Valid_o(decodedPacketValid[1]), 
        .decodedPacket1_o({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, \decodedPacket[1][120] , 
        \decodedPacket[1][119] , \decodedPacket[1][118] , 
        SYNOPSYS_UNCONNECTED__9, \decodedPacket[1][116] , 
        \decodedPacket[1][115] , \decodedPacket[1][114] , 
        \decodedPacket[1][113] , \decodedPacket[1][112] , 
        \decodedPacket[1][111] , \decodedPacket[1][110] , 
        \decodedPacket[1][109] , \decodedPacket[1][108] , 
        \decodedPacket[1][107] , \decodedPacket[1][106] , 
        \decodedPacket[1][105] , \decodedPacket[1][104] , 
        \decodedPacket[1][103] , \decodedPacket[1][102] , 
        \decodedPacket[1][101] , \decodedPacket[1][100] , 
        \decodedPacket[1][99] , \decodedPacket[1][98] , \decodedPacket[1][97] , 
        \decodedPacket[1][96] , \decodedPacket[1][95] , \decodedPacket[1][94] , 
        \decodedPacket[1][93] , \decodedPacket[1][92] , \decodedPacket[1][91] , 
        \decodedPacket[1][90] , \decodedPacket[1][89] , \decodedPacket[1][88] , 
        \decodedPacket[1][87] , \decodedPacket[1][86] , \decodedPacket[1][85] , 
        \decodedPacket[1][84] , \decodedPacket[1][83] , \decodedPacket[1][82] , 
        \decodedPacket[1][81] , \decodedPacket[1][80] , \decodedPacket[1][79] , 
        \decodedPacket[1][78] , \decodedPacket[1][77] , \decodedPacket[1][76] , 
        \decodedPacket[1][75] , \decodedPacket[1][74] , \decodedPacket[1][73] , 
        \decodedPacket[1][72] , \decodedPacket[1][71] , \decodedPacket[1][70] , 
        \decodedPacket[1][69] , \decodedPacket[1][68] , \decodedPacket[1][67] , 
        \decodedPacket[1][66] , \decodedPacket[1][65] , \decodedPacket[1][64] , 
        \decodedPacket[1][63] , \decodedPacket[1][62] , \decodedPacket[1][61] , 
        \decodedPacket[1][60] , \decodedPacket[1][59] , \decodedPacket[1][58] , 
        \decodedPacket[1][57] , \decodedPacket[1][56] , \decodedPacket[1][55] , 
        \decodedPacket[1][54] , \decodedPacket[1][53] , \decodedPacket[1][52] , 
        \decodedPacket[1][51] , \decodedPacket[1][50] , \decodedPacket[1][49] , 
        \decodedPacket[1][48] , \decodedPacket[1][47] , \decodedPacket[1][46] , 
        \decodedPacket[1][45] , \decodedPacket[1][44] , \decodedPacket[1][43] , 
        \decodedPacket[1][42] , \decodedPacket[1][41] , \decodedPacket[1][40] , 
        \decodedPacket[1][39] , \decodedPacket[1][38] , \decodedPacket[1][37] , 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        \decodedPacket[1][4] , \decodedPacket[1][3] , \decodedPacket[1][2] , 
        \decodedPacket[1][1] , \decodedPacket[1][0] }) );
  Decode_PISA_3 decode1_PISA ( .instPacketValid_i(inst1PacketValid_i), 
        .instPacket_i(inst1Packet_i), .decodedPacket0Valid_o(
        decodedPacketValid[2]), .decodedPacket0_o({SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, \decodedPacket[2][121] , 
        \decodedPacket[2][120] , \decodedPacket[2][119] , 
        \decodedPacket[2][118] , \decodedPacket[2][117] , 
        \decodedPacket[2][116] , \decodedPacket[2][115] , 
        \decodedPacket[2][114] , \decodedPacket[2][113] , 
        \decodedPacket[2][112] , \decodedPacket[2][111] , 
        \decodedPacket[2][110] , \decodedPacket[2][109] , 
        \decodedPacket[2][108] , \decodedPacket[2][107] , 
        \decodedPacket[2][106] , \decodedPacket[2][105] , 
        \decodedPacket[2][104] , \decodedPacket[2][103] , 
        \decodedPacket[2][102] , \decodedPacket[2][101] , 
        \decodedPacket[2][100] , \decodedPacket[2][99] , 
        \decodedPacket[2][98] , \decodedPacket[2][97] , \decodedPacket[2][96] , 
        \decodedPacket[2][95] , \decodedPacket[2][94] , \decodedPacket[2][93] , 
        \decodedPacket[2][92] , \decodedPacket[2][91] , \decodedPacket[2][90] , 
        \decodedPacket[2][89] , \decodedPacket[2][88] , \decodedPacket[2][87] , 
        \decodedPacket[2][86] , \decodedPacket[2][85] , \decodedPacket[2][84] , 
        \decodedPacket[2][83] , \decodedPacket[2][82] , \decodedPacket[2][81] , 
        \decodedPacket[2][80] , \decodedPacket[2][79] , \decodedPacket[2][78] , 
        \decodedPacket[2][77] , \decodedPacket[2][76] , \decodedPacket[2][75] , 
        \decodedPacket[2][74] , \decodedPacket[2][73] , \decodedPacket[2][72] , 
        \decodedPacket[2][71] , \decodedPacket[2][70] , \decodedPacket[2][69] , 
        \decodedPacket[2][68] , \decodedPacket[2][67] , \decodedPacket[2][66] , 
        \decodedPacket[2][65] , \decodedPacket[2][64] , \decodedPacket[2][63] , 
        \decodedPacket[2][62] , \decodedPacket[2][61] , \decodedPacket[2][60] , 
        \decodedPacket[2][59] , \decodedPacket[2][58] , \decodedPacket[2][57] , 
        \decodedPacket[2][56] , \decodedPacket[2][55] , \decodedPacket[2][54] , 
        \decodedPacket[2][53] , \decodedPacket[2][52] , \decodedPacket[2][51] , 
        \decodedPacket[2][50] , \decodedPacket[2][49] , \decodedPacket[2][48] , 
        \decodedPacket[2][47] , \decodedPacket[2][46] , \decodedPacket[2][45] , 
        \decodedPacket[2][44] , \decodedPacket[2][43] , \decodedPacket[2][42] , 
        \decodedPacket[2][41] , \decodedPacket[2][40] , \decodedPacket[2][39] , 
        \decodedPacket[2][38] , \decodedPacket[2][37] , \decodedPacket[2][36] , 
        \decodedPacket[2][35] , \decodedPacket[2][34] , \decodedPacket[2][33] , 
        \decodedPacket[2][32] , \decodedPacket[2][31] , \decodedPacket[2][30] , 
        \decodedPacket[2][29] , \decodedPacket[2][28] , \decodedPacket[2][27] , 
        \decodedPacket[2][26] , \decodedPacket[2][25] , \decodedPacket[2][24] , 
        \decodedPacket[2][23] , \decodedPacket[2][22] , \decodedPacket[2][21] , 
        \decodedPacket[2][20] , \decodedPacket[2][19] , \decodedPacket[2][18] , 
        \decodedPacket[2][17] , \decodedPacket[2][16] , \decodedPacket[2][15] , 
        \decodedPacket[2][14] , \decodedPacket[2][13] , \decodedPacket[2][12] , 
        \decodedPacket[2][11] , \decodedPacket[2][10] , \decodedPacket[2][9] , 
        \decodedPacket[2][8] , \decodedPacket[2][7] , \decodedPacket[2][6] , 
        \decodedPacket[2][5] , \decodedPacket[2][4] , \decodedPacket[2][3] , 
        \decodedPacket[2][2] , \decodedPacket[2][1] , \decodedPacket[2][0] }), 
        .decodedPacket1Valid_o(decodedPacketValid[3]), .decodedPacket1_o({
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, \decodedPacket[3][120] , 
        \decodedPacket[3][119] , \decodedPacket[3][118] , 
        SYNOPSYS_UNCONNECTED__51, \decodedPacket[3][116] , 
        \decodedPacket[3][115] , \decodedPacket[3][114] , 
        \decodedPacket[3][113] , \decodedPacket[3][112] , 
        \decodedPacket[3][111] , \decodedPacket[3][110] , 
        \decodedPacket[3][109] , \decodedPacket[3][108] , 
        \decodedPacket[3][107] , \decodedPacket[3][106] , 
        \decodedPacket[3][105] , \decodedPacket[3][104] , 
        \decodedPacket[3][103] , \decodedPacket[3][102] , 
        \decodedPacket[3][101] , \decodedPacket[3][100] , 
        \decodedPacket[3][99] , \decodedPacket[3][98] , \decodedPacket[3][97] , 
        \decodedPacket[3][96] , \decodedPacket[3][95] , \decodedPacket[3][94] , 
        \decodedPacket[3][93] , \decodedPacket[3][92] , \decodedPacket[3][91] , 
        \decodedPacket[3][90] , \decodedPacket[3][89] , \decodedPacket[3][88] , 
        \decodedPacket[3][87] , \decodedPacket[3][86] , \decodedPacket[3][85] , 
        \decodedPacket[3][84] , \decodedPacket[3][83] , \decodedPacket[3][82] , 
        \decodedPacket[3][81] , \decodedPacket[3][80] , \decodedPacket[3][79] , 
        \decodedPacket[3][78] , \decodedPacket[3][77] , \decodedPacket[3][76] , 
        \decodedPacket[3][75] , \decodedPacket[3][74] , \decodedPacket[3][73] , 
        \decodedPacket[3][72] , \decodedPacket[3][71] , \decodedPacket[3][70] , 
        \decodedPacket[3][69] , \decodedPacket[3][68] , \decodedPacket[3][67] , 
        \decodedPacket[3][66] , \decodedPacket[3][65] , \decodedPacket[3][64] , 
        \decodedPacket[3][63] , \decodedPacket[3][62] , \decodedPacket[3][61] , 
        \decodedPacket[3][60] , \decodedPacket[3][59] , \decodedPacket[3][58] , 
        \decodedPacket[3][57] , \decodedPacket[3][56] , \decodedPacket[3][55] , 
        \decodedPacket[3][54] , \decodedPacket[3][53] , \decodedPacket[3][52] , 
        \decodedPacket[3][51] , \decodedPacket[3][50] , \decodedPacket[3][49] , 
        \decodedPacket[3][48] , \decodedPacket[3][47] , \decodedPacket[3][46] , 
        \decodedPacket[3][45] , \decodedPacket[3][44] , \decodedPacket[3][43] , 
        \decodedPacket[3][42] , \decodedPacket[3][41] , \decodedPacket[3][40] , 
        \decodedPacket[3][39] , \decodedPacket[3][38] , \decodedPacket[3][37] , 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        \decodedPacket[3][4] , \decodedPacket[3][3] , \decodedPacket[3][2] , 
        \decodedPacket[3][1] , \decodedPacket[3][0] }) );
  Decode_PISA_2 decode2_PISA ( .instPacketValid_i(inst2PacketValid_i), 
        .instPacket_i(inst2Packet_i), .decodedPacket0Valid_o(
        decodedPacketValid[4]), .decodedPacket0_o({SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, \decodedPacket[4][121] , 
        \decodedPacket[4][120] , \decodedPacket[4][119] , 
        \decodedPacket[4][118] , \decodedPacket[4][117] , 
        \decodedPacket[4][116] , \decodedPacket[4][115] , 
        \decodedPacket[4][114] , \decodedPacket[4][113] , 
        \decodedPacket[4][112] , \decodedPacket[4][111] , 
        \decodedPacket[4][110] , \decodedPacket[4][109] , 
        \decodedPacket[4][108] , \decodedPacket[4][107] , 
        \decodedPacket[4][106] , \decodedPacket[4][105] , 
        \decodedPacket[4][104] , \decodedPacket[4][103] , 
        \decodedPacket[4][102] , \decodedPacket[4][101] , 
        \decodedPacket[4][100] , \decodedPacket[4][99] , 
        \decodedPacket[4][98] , \decodedPacket[4][97] , \decodedPacket[4][96] , 
        \decodedPacket[4][95] , \decodedPacket[4][94] , \decodedPacket[4][93] , 
        \decodedPacket[4][92] , \decodedPacket[4][91] , \decodedPacket[4][90] , 
        \decodedPacket[4][89] , \decodedPacket[4][88] , \decodedPacket[4][87] , 
        \decodedPacket[4][86] , \decodedPacket[4][85] , \decodedPacket[4][84] , 
        \decodedPacket[4][83] , \decodedPacket[4][82] , \decodedPacket[4][81] , 
        \decodedPacket[4][80] , \decodedPacket[4][79] , \decodedPacket[4][78] , 
        \decodedPacket[4][77] , \decodedPacket[4][76] , \decodedPacket[4][75] , 
        \decodedPacket[4][74] , \decodedPacket[4][73] , \decodedPacket[4][72] , 
        \decodedPacket[4][71] , \decodedPacket[4][70] , \decodedPacket[4][69] , 
        \decodedPacket[4][68] , \decodedPacket[4][67] , \decodedPacket[4][66] , 
        \decodedPacket[4][65] , \decodedPacket[4][64] , \decodedPacket[4][63] , 
        \decodedPacket[4][62] , \decodedPacket[4][61] , \decodedPacket[4][60] , 
        \decodedPacket[4][59] , \decodedPacket[4][58] , \decodedPacket[4][57] , 
        \decodedPacket[4][56] , \decodedPacket[4][55] , \decodedPacket[4][54] , 
        \decodedPacket[4][53] , \decodedPacket[4][52] , \decodedPacket[4][51] , 
        \decodedPacket[4][50] , \decodedPacket[4][49] , \decodedPacket[4][48] , 
        \decodedPacket[4][47] , \decodedPacket[4][46] , \decodedPacket[4][45] , 
        \decodedPacket[4][44] , \decodedPacket[4][43] , \decodedPacket[4][42] , 
        \decodedPacket[4][41] , \decodedPacket[4][40] , \decodedPacket[4][39] , 
        \decodedPacket[4][38] , \decodedPacket[4][37] , \decodedPacket[4][36] , 
        \decodedPacket[4][35] , \decodedPacket[4][34] , \decodedPacket[4][33] , 
        \decodedPacket[4][32] , \decodedPacket[4][31] , \decodedPacket[4][30] , 
        \decodedPacket[4][29] , \decodedPacket[4][28] , \decodedPacket[4][27] , 
        \decodedPacket[4][26] , \decodedPacket[4][25] , \decodedPacket[4][24] , 
        \decodedPacket[4][23] , \decodedPacket[4][22] , \decodedPacket[4][21] , 
        \decodedPacket[4][20] , \decodedPacket[4][19] , \decodedPacket[4][18] , 
        \decodedPacket[4][17] , \decodedPacket[4][16] , \decodedPacket[4][15] , 
        \decodedPacket[4][14] , \decodedPacket[4][13] , \decodedPacket[4][12] , 
        \decodedPacket[4][11] , \decodedPacket[4][10] , \decodedPacket[4][9] , 
        \decodedPacket[4][8] , \decodedPacket[4][7] , \decodedPacket[4][6] , 
        \decodedPacket[4][5] , \decodedPacket[4][4] , \decodedPacket[4][3] , 
        \decodedPacket[4][2] , \decodedPacket[4][1] , \decodedPacket[4][0] }), 
        .decodedPacket1Valid_o(decodedPacketValid[5]), .decodedPacket1_o({
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, \decodedPacket[5][120] , 
        \decodedPacket[5][119] , \decodedPacket[5][118] , 
        SYNOPSYS_UNCONNECTED__93, \decodedPacket[5][116] , 
        \decodedPacket[5][115] , \decodedPacket[5][114] , 
        \decodedPacket[5][113] , \decodedPacket[5][112] , 
        \decodedPacket[5][111] , \decodedPacket[5][110] , 
        \decodedPacket[5][109] , \decodedPacket[5][108] , 
        \decodedPacket[5][107] , \decodedPacket[5][106] , 
        \decodedPacket[5][105] , \decodedPacket[5][104] , 
        \decodedPacket[5][103] , \decodedPacket[5][102] , 
        \decodedPacket[5][101] , \decodedPacket[5][100] , 
        \decodedPacket[5][99] , \decodedPacket[5][98] , \decodedPacket[5][97] , 
        \decodedPacket[5][96] , \decodedPacket[5][95] , \decodedPacket[5][94] , 
        \decodedPacket[5][93] , \decodedPacket[5][92] , \decodedPacket[5][91] , 
        \decodedPacket[5][90] , \decodedPacket[5][89] , \decodedPacket[5][88] , 
        \decodedPacket[5][87] , \decodedPacket[5][86] , \decodedPacket[5][85] , 
        \decodedPacket[5][84] , \decodedPacket[5][83] , \decodedPacket[5][82] , 
        \decodedPacket[5][81] , \decodedPacket[5][80] , \decodedPacket[5][79] , 
        \decodedPacket[5][78] , \decodedPacket[5][77] , \decodedPacket[5][76] , 
        \decodedPacket[5][75] , \decodedPacket[5][74] , \decodedPacket[5][73] , 
        \decodedPacket[5][72] , \decodedPacket[5][71] , \decodedPacket[5][70] , 
        \decodedPacket[5][69] , \decodedPacket[5][68] , \decodedPacket[5][67] , 
        \decodedPacket[5][66] , \decodedPacket[5][65] , \decodedPacket[5][64] , 
        \decodedPacket[5][63] , \decodedPacket[5][62] , \decodedPacket[5][61] , 
        \decodedPacket[5][60] , \decodedPacket[5][59] , \decodedPacket[5][58] , 
        \decodedPacket[5][57] , \decodedPacket[5][56] , \decodedPacket[5][55] , 
        \decodedPacket[5][54] , \decodedPacket[5][53] , \decodedPacket[5][52] , 
        \decodedPacket[5][51] , \decodedPacket[5][50] , \decodedPacket[5][49] , 
        \decodedPacket[5][48] , \decodedPacket[5][47] , \decodedPacket[5][46] , 
        \decodedPacket[5][45] , \decodedPacket[5][44] , \decodedPacket[5][43] , 
        \decodedPacket[5][42] , \decodedPacket[5][41] , \decodedPacket[5][40] , 
        \decodedPacket[5][39] , \decodedPacket[5][38] , \decodedPacket[5][37] , 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        \decodedPacket[5][4] , \decodedPacket[5][3] , \decodedPacket[5][2] , 
        \decodedPacket[5][1] , \decodedPacket[5][0] }) );
  Decode_PISA_1 decode3_PISA ( .instPacketValid_i(inst3PacketValid_i), 
        .instPacket_i(inst3Packet_i), .decodedPacket0Valid_o(
        decodedPacketValid[6]), .decodedPacket0_o({SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, \decodedPacket[6][121] , 
        \decodedPacket[6][120] , \decodedPacket[6][119] , 
        \decodedPacket[6][118] , \decodedPacket[6][117] , 
        \decodedPacket[6][116] , \decodedPacket[6][115] , 
        \decodedPacket[6][114] , \decodedPacket[6][113] , 
        \decodedPacket[6][112] , \decodedPacket[6][111] , 
        \decodedPacket[6][110] , \decodedPacket[6][109] , 
        \decodedPacket[6][108] , \decodedPacket[6][107] , 
        \decodedPacket[6][106] , \decodedPacket[6][105] , 
        \decodedPacket[6][104] , \decodedPacket[6][103] , 
        \decodedPacket[6][102] , \decodedPacket[6][101] , 
        \decodedPacket[6][100] , \decodedPacket[6][99] , 
        \decodedPacket[6][98] , \decodedPacket[6][97] , \decodedPacket[6][96] , 
        \decodedPacket[6][95] , \decodedPacket[6][94] , \decodedPacket[6][93] , 
        \decodedPacket[6][92] , \decodedPacket[6][91] , \decodedPacket[6][90] , 
        \decodedPacket[6][89] , \decodedPacket[6][88] , \decodedPacket[6][87] , 
        \decodedPacket[6][86] , \decodedPacket[6][85] , \decodedPacket[6][84] , 
        \decodedPacket[6][83] , \decodedPacket[6][82] , \decodedPacket[6][81] , 
        \decodedPacket[6][80] , \decodedPacket[6][79] , \decodedPacket[6][78] , 
        \decodedPacket[6][77] , \decodedPacket[6][76] , \decodedPacket[6][75] , 
        \decodedPacket[6][74] , \decodedPacket[6][73] , \decodedPacket[6][72] , 
        \decodedPacket[6][71] , \decodedPacket[6][70] , \decodedPacket[6][69] , 
        \decodedPacket[6][68] , \decodedPacket[6][67] , \decodedPacket[6][66] , 
        \decodedPacket[6][65] , \decodedPacket[6][64] , \decodedPacket[6][63] , 
        \decodedPacket[6][62] , \decodedPacket[6][61] , \decodedPacket[6][60] , 
        \decodedPacket[6][59] , \decodedPacket[6][58] , \decodedPacket[6][57] , 
        \decodedPacket[6][56] , \decodedPacket[6][55] , \decodedPacket[6][54] , 
        \decodedPacket[6][53] , \decodedPacket[6][52] , \decodedPacket[6][51] , 
        \decodedPacket[6][50] , \decodedPacket[6][49] , \decodedPacket[6][48] , 
        \decodedPacket[6][47] , \decodedPacket[6][46] , \decodedPacket[6][45] , 
        \decodedPacket[6][44] , \decodedPacket[6][43] , \decodedPacket[6][42] , 
        \decodedPacket[6][41] , \decodedPacket[6][40] , \decodedPacket[6][39] , 
        \decodedPacket[6][38] , \decodedPacket[6][37] , \decodedPacket[6][36] , 
        \decodedPacket[6][35] , \decodedPacket[6][34] , \decodedPacket[6][33] , 
        \decodedPacket[6][32] , \decodedPacket[6][31] , \decodedPacket[6][30] , 
        \decodedPacket[6][29] , \decodedPacket[6][28] , \decodedPacket[6][27] , 
        \decodedPacket[6][26] , \decodedPacket[6][25] , \decodedPacket[6][24] , 
        \decodedPacket[6][23] , \decodedPacket[6][22] , \decodedPacket[6][21] , 
        \decodedPacket[6][20] , \decodedPacket[6][19] , \decodedPacket[6][18] , 
        \decodedPacket[6][17] , \decodedPacket[6][16] , \decodedPacket[6][15] , 
        \decodedPacket[6][14] , \decodedPacket[6][13] , \decodedPacket[6][12] , 
        \decodedPacket[6][11] , \decodedPacket[6][10] , \decodedPacket[6][9] , 
        \decodedPacket[6][8] , \decodedPacket[6][7] , \decodedPacket[6][6] , 
        \decodedPacket[6][5] , \decodedPacket[6][4] , \decodedPacket[6][3] , 
        \decodedPacket[6][2] , \decodedPacket[6][1] , \decodedPacket[6][0] }), 
        .decodedPacket1Valid_o(decodedPacketValid[7]), .decodedPacket1_o({
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, \decodedPacket[7][120] , 
        \decodedPacket[7][119] , \decodedPacket[7][118] , 
        SYNOPSYS_UNCONNECTED__135, \decodedPacket[7][116] , 
        \decodedPacket[7][115] , \decodedPacket[7][114] , 
        \decodedPacket[7][113] , \decodedPacket[7][112] , 
        \decodedPacket[7][111] , \decodedPacket[7][110] , 
        \decodedPacket[7][109] , \decodedPacket[7][108] , 
        \decodedPacket[7][107] , \decodedPacket[7][106] , 
        \decodedPacket[7][105] , \decodedPacket[7][104] , 
        \decodedPacket[7][103] , \decodedPacket[7][102] , 
        \decodedPacket[7][101] , \decodedPacket[7][100] , 
        \decodedPacket[7][99] , \decodedPacket[7][98] , \decodedPacket[7][97] , 
        \decodedPacket[7][96] , \decodedPacket[7][95] , \decodedPacket[7][94] , 
        \decodedPacket[7][93] , \decodedPacket[7][92] , \decodedPacket[7][91] , 
        \decodedPacket[7][90] , \decodedPacket[7][89] , \decodedPacket[7][88] , 
        \decodedPacket[7][87] , \decodedPacket[7][86] , \decodedPacket[7][85] , 
        \decodedPacket[7][84] , \decodedPacket[7][83] , \decodedPacket[7][82] , 
        \decodedPacket[7][81] , \decodedPacket[7][80] , \decodedPacket[7][79] , 
        \decodedPacket[7][78] , \decodedPacket[7][77] , \decodedPacket[7][76] , 
        \decodedPacket[7][75] , \decodedPacket[7][74] , \decodedPacket[7][73] , 
        \decodedPacket[7][72] , \decodedPacket[7][71] , \decodedPacket[7][70] , 
        \decodedPacket[7][69] , \decodedPacket[7][68] , \decodedPacket[7][67] , 
        \decodedPacket[7][66] , \decodedPacket[7][65] , \decodedPacket[7][64] , 
        \decodedPacket[7][63] , \decodedPacket[7][62] , \decodedPacket[7][61] , 
        \decodedPacket[7][60] , \decodedPacket[7][59] , \decodedPacket[7][58] , 
        \decodedPacket[7][57] , \decodedPacket[7][56] , \decodedPacket[7][55] , 
        \decodedPacket[7][54] , \decodedPacket[7][53] , \decodedPacket[7][52] , 
        \decodedPacket[7][51] , \decodedPacket[7][50] , \decodedPacket[7][49] , 
        \decodedPacket[7][48] , \decodedPacket[7][47] , \decodedPacket[7][46] , 
        \decodedPacket[7][45] , \decodedPacket[7][44] , \decodedPacket[7][43] , 
        \decodedPacket[7][42] , \decodedPacket[7][41] , \decodedPacket[7][40] , 
        \decodedPacket[7][39] , \decodedPacket[7][38] , \decodedPacket[7][37] , 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        \decodedPacket[7][4] , \decodedPacket[7][3] , \decodedPacket[7][2] , 
        \decodedPacket[7][1] , \decodedPacket[7][0] }) );
  INVX0 U5859 ( .INP(1'b1), .ZN(decodedPacket7_o[122]) );
  INVX0 U5861 ( .INP(1'b1), .ZN(decodedPacket7_o[123]) );
  INVX0 U5863 ( .INP(1'b1), .ZN(decodedPacket7_o[124]) );
  INVX0 U5865 ( .INP(1'b1), .ZN(decodedPacket7_o[125]) );
  INVX0 U5867 ( .INP(1'b1), .ZN(decodedPacket6_o[122]) );
  INVX0 U5869 ( .INP(1'b1), .ZN(decodedPacket6_o[123]) );
  INVX0 U5871 ( .INP(1'b1), .ZN(decodedPacket6_o[124]) );
  INVX0 U5873 ( .INP(1'b1), .ZN(decodedPacket6_o[125]) );
  INVX0 U5875 ( .INP(1'b1), .ZN(decodedPacket5_o[122]) );
  INVX0 U5877 ( .INP(1'b1), .ZN(decodedPacket5_o[123]) );
  INVX0 U5879 ( .INP(1'b1), .ZN(decodedPacket5_o[124]) );
  INVX0 U5881 ( .INP(1'b1), .ZN(decodedPacket5_o[125]) );
  INVX0 U5883 ( .INP(1'b1), .ZN(decodedPacket4_o[122]) );
  INVX0 U5885 ( .INP(1'b1), .ZN(decodedPacket4_o[123]) );
  INVX0 U5887 ( .INP(1'b1), .ZN(decodedPacket4_o[124]) );
  INVX0 U5889 ( .INP(1'b1), .ZN(decodedPacket4_o[125]) );
  INVX0 U5891 ( .INP(1'b1), .ZN(decodedPacket3_o[122]) );
  INVX0 U5893 ( .INP(1'b1), .ZN(decodedPacket3_o[123]) );
  INVX0 U5895 ( .INP(1'b1), .ZN(decodedPacket3_o[124]) );
  INVX0 U5897 ( .INP(1'b1), .ZN(decodedPacket3_o[125]) );
  INVX0 U5899 ( .INP(1'b1), .ZN(decodedPacket2_o[122]) );
  INVX0 U5901 ( .INP(1'b1), .ZN(decodedPacket2_o[123]) );
  INVX0 U5903 ( .INP(1'b1), .ZN(decodedPacket2_o[124]) );
  INVX0 U5905 ( .INP(1'b1), .ZN(decodedPacket2_o[125]) );
  INVX0 U5907 ( .INP(1'b1), .ZN(decodedPacket1_o[122]) );
  INVX0 U5909 ( .INP(1'b1), .ZN(decodedPacket1_o[123]) );
  INVX0 U5911 ( .INP(1'b1), .ZN(decodedPacket1_o[124]) );
  INVX0 U5913 ( .INP(1'b1), .ZN(decodedPacket1_o[125]) );
  INVX0 U5915 ( .INP(1'b1), .ZN(decodedPacket0_o[122]) );
  INVX0 U5917 ( .INP(1'b1), .ZN(decodedPacket0_o[123]) );
  INVX0 U5919 ( .INP(1'b1), .ZN(decodedPacket0_o[124]) );
  INVX0 U5921 ( .INP(1'b1), .ZN(decodedPacket0_o[125]) );
  AND4X1 U5923 ( .IN1(n1754), .IN2(decodedPacketValid[4]), .IN3(N2172), .IN4(
        n5990), .Q(n4910) );
  NAND2X1 U5924 ( .IN1(n4837), .IN2(n5192), .QN(n4066) );
  INVX0 U5925 ( .INP(\decodedPacket[3][114] ), .ZN(n5937) );
  INVX0 U5926 ( .INP(\decodedPacket[5][114] ), .ZN(n5952) );
  INVX0 U5927 ( .INP(\decodedPacket[7][114] ), .ZN(n5967) );
  INVX0 U5928 ( .INP(\decodedPacket[4][118] ), .ZN(n6220) );
  INVX0 U5929 ( .INP(\decodedPacket[6][118] ), .ZN(n6374) );
  AND4X1 U5930 ( .IN1(decodedPacketValid[5]), .IN2(n2907), .IN3(n5994), .IN4(
        n5989), .Q(n4911) );
  AND4X1 U5931 ( .IN1(decodedPacketValid[5]), .IN2(N4308), .IN3(n2907), .IN4(
        n5989), .Q(n4912) );
  AND4X1 U5932 ( .IN1(decodedPacketValid[5]), .IN2(N4309), .IN3(n2907), .IN4(
        n5994), .Q(n4913) );
  AND4X1 U5933 ( .IN1(decodedPacketValid[5]), .IN2(N4309), .IN3(N4308), .IN4(
        n2907), .Q(n4914) );
  AND4X1 U5934 ( .IN1(n1755), .IN2(decodedPacketValid[5]), .IN3(N4308), .IN4(
        n5989), .Q(n4915) );
  AND4X1 U5935 ( .IN1(n1755), .IN2(decodedPacketValid[5]), .IN3(N4309), .IN4(
        N4308), .Q(n4916) );
  AND4X1 U5936 ( .IN1(n1755), .IN2(decodedPacketValid[5]), .IN3(n5994), .IN4(
        n5989), .Q(n4917) );
  AND4X1 U5937 ( .IN1(n1755), .IN2(decodedPacketValid[5]), .IN3(N4309), .IN4(
        n5994), .Q(n4918) );
  AND4X1 U5938 ( .IN1(n5986), .IN2(decodedPacketValid[3]), .IN3(N1069), .IN4(
        n5996), .Q(n4919) );
  AND2X1 U5939 ( .IN1(\decodedPacket[4][11] ), .IN2(n5529), .Q(n4920) );
  AND2X1 U5940 ( .IN1(\decodedPacket[4][13] ), .IN2(n5529), .Q(n4921) );
  AND2X1 U5941 ( .IN1(\decodedPacket[4][14] ), .IN2(n5529), .Q(n4922) );
  AND2X1 U5942 ( .IN1(\decodedPacket[4][15] ), .IN2(n5529), .Q(n4923) );
  AND2X1 U5943 ( .IN1(\decodedPacket[4][16] ), .IN2(n5529), .Q(n4924) );
  AND2X1 U5944 ( .IN1(\decodedPacket[4][17] ), .IN2(n5529), .Q(n4925) );
  AND2X1 U5945 ( .IN1(\decodedPacket[4][18] ), .IN2(n5529), .Q(n4926) );
  AND2X1 U5946 ( .IN1(\decodedPacket[4][19] ), .IN2(n5529), .Q(n4927) );
  AND2X1 U5947 ( .IN1(\decodedPacket[4][20] ), .IN2(n5529), .Q(n4928) );
  AND2X1 U5948 ( .IN1(\decodedPacket[4][21] ), .IN2(n5529), .Q(n4929) );
  AND2X1 U5949 ( .IN1(\decodedPacket[4][23] ), .IN2(n5529), .Q(n4930) );
  AND2X1 U5950 ( .IN1(\decodedPacket[4][24] ), .IN2(n5529), .Q(n4931) );
  AND2X1 U5951 ( .IN1(\decodedPacket[4][26] ), .IN2(n5529), .Q(n4932) );
  AND2X1 U5952 ( .IN1(\decodedPacket[4][117] ), .IN2(n5528), .Q(n4933) );
  AND2X1 U5953 ( .IN1(\decodedPacket[4][27] ), .IN2(n5528), .Q(n4934) );
  AND2X1 U5954 ( .IN1(\decodedPacket[4][28] ), .IN2(n5528), .Q(n4935) );
  AND2X1 U5955 ( .IN1(\decodedPacket[4][29] ), .IN2(n5528), .Q(n4936) );
  AND2X1 U5956 ( .IN1(\decodedPacket[4][30] ), .IN2(n5528), .Q(n4937) );
  AND2X1 U5957 ( .IN1(\decodedPacket[4][31] ), .IN2(n5528), .Q(n4938) );
  AND2X1 U5958 ( .IN1(\decodedPacket[4][32] ), .IN2(n5528), .Q(n4939) );
  AND2X1 U5959 ( .IN1(\decodedPacket[4][33] ), .IN2(n5528), .Q(n4940) );
  AND2X1 U5960 ( .IN1(\decodedPacket[4][34] ), .IN2(n5528), .Q(n4941) );
  AND2X1 U5961 ( .IN1(\decodedPacket[4][35] ), .IN2(n5528), .Q(n4942) );
  AND2X1 U5962 ( .IN1(\decodedPacket[4][36] ), .IN2(n5528), .Q(n4943) );
  AND2X1 U5963 ( .IN1(\decodedPacket[4][25] ), .IN2(n5528), .Q(n4944) );
  AND2X1 U5964 ( .IN1(\decodedPacket[4][11] ), .IN2(n5352), .Q(n4945) );
  AND2X1 U5965 ( .IN1(\decodedPacket[4][13] ), .IN2(n5352), .Q(n4946) );
  AND2X1 U5966 ( .IN1(\decodedPacket[4][14] ), .IN2(n5352), .Q(n4947) );
  AND2X1 U5967 ( .IN1(\decodedPacket[4][11] ), .IN2(n5411), .Q(n4948) );
  AND2X1 U5968 ( .IN1(\decodedPacket[4][13] ), .IN2(n5411), .Q(n4949) );
  AND2X1 U5969 ( .IN1(\decodedPacket[4][14] ), .IN2(n5411), .Q(n4950) );
  AND2X1 U5970 ( .IN1(\decodedPacket[4][11] ), .IN2(n5470), .Q(n4951) );
  AND2X1 U5971 ( .IN1(\decodedPacket[4][13] ), .IN2(n5470), .Q(n4952) );
  AND2X1 U5972 ( .IN1(\decodedPacket[4][14] ), .IN2(n5470), .Q(n4953) );
  AND2X1 U5973 ( .IN1(\decodedPacket[4][15] ), .IN2(n5352), .Q(n4954) );
  AND2X1 U5974 ( .IN1(\decodedPacket[4][16] ), .IN2(n5352), .Q(n4955) );
  AND2X1 U5975 ( .IN1(\decodedPacket[4][17] ), .IN2(n5352), .Q(n4956) );
  AND2X1 U5976 ( .IN1(\decodedPacket[4][18] ), .IN2(n5352), .Q(n4957) );
  AND2X1 U5977 ( .IN1(\decodedPacket[4][19] ), .IN2(n5352), .Q(n4958) );
  AND2X1 U5978 ( .IN1(\decodedPacket[4][20] ), .IN2(n5352), .Q(n4959) );
  AND2X1 U5979 ( .IN1(\decodedPacket[4][21] ), .IN2(n5352), .Q(n4960) );
  AND2X1 U5980 ( .IN1(\decodedPacket[4][22] ), .IN2(n5352), .Q(n4961) );
  AND2X1 U5981 ( .IN1(\decodedPacket[4][23] ), .IN2(n5352), .Q(n4962) );
  AND2X1 U5982 ( .IN1(\decodedPacket[4][24] ), .IN2(n5352), .Q(n4963) );
  AND2X1 U5983 ( .IN1(\decodedPacket[4][26] ), .IN2(n5352), .Q(n4964) );
  AND2X1 U5984 ( .IN1(\decodedPacket[4][15] ), .IN2(n5411), .Q(n4965) );
  AND2X1 U5985 ( .IN1(\decodedPacket[4][16] ), .IN2(n5411), .Q(n4966) );
  AND2X1 U5986 ( .IN1(\decodedPacket[4][17] ), .IN2(n5411), .Q(n4967) );
  AND2X1 U5987 ( .IN1(\decodedPacket[4][18] ), .IN2(n5411), .Q(n4968) );
  AND2X1 U5988 ( .IN1(\decodedPacket[4][19] ), .IN2(n5411), .Q(n4969) );
  AND2X1 U5989 ( .IN1(\decodedPacket[4][20] ), .IN2(n5411), .Q(n4970) );
  AND2X1 U5990 ( .IN1(\decodedPacket[4][21] ), .IN2(n5411), .Q(n4971) );
  AND2X1 U5991 ( .IN1(\decodedPacket[4][22] ), .IN2(n5411), .Q(n4972) );
  AND2X1 U5992 ( .IN1(\decodedPacket[4][23] ), .IN2(n5411), .Q(n4973) );
  AND2X1 U5993 ( .IN1(\decodedPacket[4][24] ), .IN2(n5411), .Q(n4974) );
  AND2X1 U5994 ( .IN1(\decodedPacket[4][26] ), .IN2(n5411), .Q(n4975) );
  AND2X1 U5995 ( .IN1(\decodedPacket[4][15] ), .IN2(n5470), .Q(n4976) );
  AND2X1 U5996 ( .IN1(\decodedPacket[4][16] ), .IN2(n5470), .Q(n4977) );
  AND2X1 U5997 ( .IN1(\decodedPacket[4][17] ), .IN2(n5470), .Q(n4978) );
  AND2X1 U5998 ( .IN1(\decodedPacket[4][18] ), .IN2(n5470), .Q(n4979) );
  AND2X1 U5999 ( .IN1(\decodedPacket[4][19] ), .IN2(n5470), .Q(n4980) );
  AND2X1 U6000 ( .IN1(\decodedPacket[4][20] ), .IN2(n5470), .Q(n4981) );
  AND2X1 U6001 ( .IN1(\decodedPacket[4][21] ), .IN2(n5470), .Q(n4982) );
  AND2X1 U6002 ( .IN1(\decodedPacket[4][22] ), .IN2(n5470), .Q(n4983) );
  AND2X1 U6003 ( .IN1(\decodedPacket[4][23] ), .IN2(n5470), .Q(n4984) );
  AND2X1 U6004 ( .IN1(\decodedPacket[4][24] ), .IN2(n5470), .Q(n4985) );
  AND2X1 U6005 ( .IN1(\decodedPacket[4][26] ), .IN2(n5470), .Q(n4986) );
  AND2X1 U6006 ( .IN1(\decodedPacket[4][22] ), .IN2(n5529), .Q(n4987) );
  AND2X1 U6007 ( .IN1(\decodedPacket[4][121] ), .IN2(n5351), .Q(n4988) );
  AND2X1 U6008 ( .IN1(\decodedPacket[4][121] ), .IN2(n5410), .Q(n4989) );
  AND2X1 U6009 ( .IN1(\decodedPacket[4][121] ), .IN2(n5469), .Q(n4990) );
  AND2X1 U6010 ( .IN1(\decodedPacket[4][121] ), .IN2(n5528), .Q(n4991) );
  AND2X1 U6011 ( .IN1(\decodedPacket[4][117] ), .IN2(n5351), .Q(n4992) );
  AND2X1 U6012 ( .IN1(\decodedPacket[4][117] ), .IN2(n5410), .Q(n4993) );
  AND2X1 U6013 ( .IN1(\decodedPacket[4][117] ), .IN2(n5469), .Q(n4994) );
  AND2X1 U6014 ( .IN1(\decodedPacket[4][27] ), .IN2(n5351), .Q(n4995) );
  AND2X1 U6015 ( .IN1(\decodedPacket[4][28] ), .IN2(n5351), .Q(n4996) );
  AND2X1 U6016 ( .IN1(\decodedPacket[4][29] ), .IN2(n5351), .Q(n4997) );
  AND2X1 U6017 ( .IN1(\decodedPacket[4][30] ), .IN2(n5351), .Q(n4998) );
  AND2X1 U6018 ( .IN1(\decodedPacket[4][31] ), .IN2(n5351), .Q(n4999) );
  AND2X1 U6019 ( .IN1(\decodedPacket[4][32] ), .IN2(n5351), .Q(n5000) );
  AND2X1 U6020 ( .IN1(\decodedPacket[4][33] ), .IN2(n5351), .Q(n5001) );
  AND2X1 U6021 ( .IN1(\decodedPacket[4][34] ), .IN2(n5351), .Q(n5002) );
  AND2X1 U6022 ( .IN1(\decodedPacket[4][35] ), .IN2(n5351), .Q(n5003) );
  AND2X1 U6023 ( .IN1(\decodedPacket[4][36] ), .IN2(n5351), .Q(n5004) );
  AND2X1 U6024 ( .IN1(\decodedPacket[4][27] ), .IN2(n5410), .Q(n5005) );
  AND2X1 U6025 ( .IN1(\decodedPacket[4][28] ), .IN2(n5410), .Q(n5006) );
  AND2X1 U6026 ( .IN1(\decodedPacket[4][29] ), .IN2(n5410), .Q(n5007) );
  AND2X1 U6027 ( .IN1(\decodedPacket[4][30] ), .IN2(n5410), .Q(n5008) );
  AND2X1 U6028 ( .IN1(\decodedPacket[4][31] ), .IN2(n5410), .Q(n5009) );
  AND2X1 U6029 ( .IN1(\decodedPacket[4][32] ), .IN2(n5410), .Q(n5010) );
  AND2X1 U6030 ( .IN1(\decodedPacket[4][33] ), .IN2(n5410), .Q(n5011) );
  AND2X1 U6031 ( .IN1(\decodedPacket[4][34] ), .IN2(n5410), .Q(n5012) );
  AND2X1 U6032 ( .IN1(\decodedPacket[4][35] ), .IN2(n5410), .Q(n5013) );
  AND2X1 U6033 ( .IN1(\decodedPacket[4][36] ), .IN2(n5410), .Q(n5014) );
  AND2X1 U6034 ( .IN1(\decodedPacket[4][27] ), .IN2(n5469), .Q(n5015) );
  AND2X1 U6035 ( .IN1(\decodedPacket[4][28] ), .IN2(n5469), .Q(n5016) );
  AND2X1 U6036 ( .IN1(\decodedPacket[4][29] ), .IN2(n5469), .Q(n5017) );
  AND2X1 U6037 ( .IN1(\decodedPacket[4][30] ), .IN2(n5469), .Q(n5018) );
  AND2X1 U6038 ( .IN1(\decodedPacket[4][31] ), .IN2(n5469), .Q(n5019) );
  AND2X1 U6039 ( .IN1(\decodedPacket[4][32] ), .IN2(n5469), .Q(n5020) );
  AND2X1 U6040 ( .IN1(\decodedPacket[4][33] ), .IN2(n5469), .Q(n5021) );
  AND2X1 U6041 ( .IN1(\decodedPacket[4][34] ), .IN2(n5469), .Q(n5022) );
  AND2X1 U6042 ( .IN1(\decodedPacket[4][35] ), .IN2(n5469), .Q(n5023) );
  AND2X1 U6043 ( .IN1(\decodedPacket[4][36] ), .IN2(n5469), .Q(n5024) );
  AND2X1 U6044 ( .IN1(\decodedPacket[4][25] ), .IN2(n5351), .Q(n5025) );
  AND2X1 U6045 ( .IN1(\decodedPacket[4][25] ), .IN2(n5410), .Q(n5026) );
  AND2X1 U6046 ( .IN1(\decodedPacket[4][25] ), .IN2(n5469), .Q(n5027) );
  OAI22X1 U6047 ( .IN1(n5626), .IN2(n2378), .IN3(n6179), .IN4(n5629), .QN(
        n5028) );
  OAI22X1 U6048 ( .IN1(n5626), .IN2(n2372), .IN3(n6178), .IN4(n5629), .QN(
        n5029) );
  OAI22X1 U6049 ( .IN1(n5626), .IN2(n2366), .IN3(n6177), .IN4(n5629), .QN(
        n5030) );
  OAI22X1 U6050 ( .IN1(n5626), .IN2(n2360), .IN3(n6176), .IN4(n5629), .QN(
        n5031) );
  OAI22X1 U6051 ( .IN1(n5626), .IN2(n2354), .IN3(n6175), .IN4(n5629), .QN(
        n5032) );
  OAI22X1 U6052 ( .IN1(n5626), .IN2(n2348), .IN3(n6174), .IN4(n5629), .QN(
        n5033) );
  OAI22X1 U6053 ( .IN1(n5626), .IN2(n2342), .IN3(n6173), .IN4(n5629), .QN(
        n5034) );
  OAI22X1 U6054 ( .IN1(n5626), .IN2(n2336), .IN3(n6172), .IN4(n5629), .QN(
        n5035) );
  OAI22X1 U6055 ( .IN1(n5626), .IN2(n2330), .IN3(n6171), .IN4(n5629), .QN(
        n5036) );
  OAI22X1 U6056 ( .IN1(n5626), .IN2(n2324), .IN3(n6170), .IN4(n5629), .QN(
        n5037) );
  OAI22X1 U6057 ( .IN1(n5626), .IN2(n2318), .IN3(n6169), .IN4(n5629), .QN(
        n5038) );
  OAI22X1 U6058 ( .IN1(n5626), .IN2(n2312), .IN3(n6168), .IN4(n5629), .QN(
        n5039) );
  OAI22X1 U6059 ( .IN1(n5626), .IN2(n2306), .IN3(n6167), .IN4(n5630), .QN(
        n5040) );
  OAI22X1 U6060 ( .IN1(n5626), .IN2(n2300), .IN3(n6166), .IN4(n5630), .QN(
        n5041) );
  OAI22X1 U6061 ( .IN1(n5624), .IN2(n1790), .IN3(n5855), .IN4(n5636), .QN(
        n5042) );
  OAI22X1 U6062 ( .IN1(n5624), .IN2(n1814), .IN3(n6217), .IN4(n5636), .QN(
        n5043) );
  OAI22X1 U6063 ( .IN1(n5627), .IN2(n2486), .IN3(n6165), .IN4(n5631), .QN(
        n5044) );
  OAI22X1 U6064 ( .IN1(n5627), .IN2(n2480), .IN3(n6164), .IN4(n5632), .QN(
        n5045) );
  OAI22X1 U6065 ( .IN1(n5627), .IN2(n2474), .IN3(n6163), .IN4(n5633), .QN(
        n5046) );
  OAI22X1 U6066 ( .IN1(n5627), .IN2(n2468), .IN3(n6162), .IN4(n5634), .QN(
        n5047) );
  OAI22X1 U6067 ( .IN1(n5627), .IN2(n2462), .IN3(n6161), .IN4(n5628), .QN(
        n5048) );
  OAI22X1 U6068 ( .IN1(n5627), .IN2(n2456), .IN3(n6192), .IN4(n5628), .QN(
        n5049) );
  OAI22X1 U6069 ( .IN1(n5627), .IN2(n2450), .IN3(n6191), .IN4(n5628), .QN(
        n5050) );
  OAI22X1 U6070 ( .IN1(n5627), .IN2(n2444), .IN3(n6190), .IN4(n5628), .QN(
        n5051) );
  OAI22X1 U6071 ( .IN1(n5627), .IN2(n2438), .IN3(n6189), .IN4(n5628), .QN(
        n5052) );
  OAI22X1 U6072 ( .IN1(n5627), .IN2(n2432), .IN3(n6188), .IN4(n5628), .QN(
        n5053) );
  OAI22X1 U6073 ( .IN1(n5627), .IN2(n2426), .IN3(n6187), .IN4(n5628), .QN(
        n5054) );
  OAI22X1 U6074 ( .IN1(n5627), .IN2(n2420), .IN3(n6186), .IN4(n5628), .QN(
        n5055) );
  OAI22X1 U6075 ( .IN1(n5627), .IN2(n2414), .IN3(n6185), .IN4(n5628), .QN(
        n5056) );
  OAI22X1 U6076 ( .IN1(n5627), .IN2(n2408), .IN3(n6184), .IN4(n5628), .QN(
        n5057) );
  OAI22X1 U6077 ( .IN1(n5627), .IN2(n2402), .IN3(n6183), .IN4(n5628), .QN(
        n5058) );
  OAI22X1 U6078 ( .IN1(n5627), .IN2(n2396), .IN3(n6182), .IN4(n5628), .QN(
        n5059) );
  OAI22X1 U6079 ( .IN1(n5627), .IN2(n2390), .IN3(n6181), .IN4(n5628), .QN(
        n5060) );
  OAI22X1 U6080 ( .IN1(n5627), .IN2(n2384), .IN3(n6180), .IN4(n5629), .QN(
        n5061) );
  OAI22X1 U6081 ( .IN1(n6190), .IN2(n5715), .IN3(n5726), .IN4(n1688), .QN(
        n5062) );
  OAI22X1 U6082 ( .IN1(n6189), .IN2(n5715), .IN3(n5726), .IN4(n1683), .QN(
        n5063) );
  OAI22X1 U6083 ( .IN1(n6188), .IN2(n5715), .IN3(n5726), .IN4(n1678), .QN(
        n5064) );
  OAI22X1 U6084 ( .IN1(n6187), .IN2(n5715), .IN3(n5726), .IN4(n1673), .QN(
        n5065) );
  OAI22X1 U6085 ( .IN1(n6186), .IN2(n5715), .IN3(n5725), .IN4(n1668), .QN(
        n5066) );
  OAI22X1 U6086 ( .IN1(n6185), .IN2(n5715), .IN3(n5725), .IN4(n1663), .QN(
        n5067) );
  OAI22X1 U6087 ( .IN1(n6184), .IN2(n5715), .IN3(n5725), .IN4(n1658), .QN(
        n5068) );
  OAI22X1 U6088 ( .IN1(n6183), .IN2(n5715), .IN3(n5725), .IN4(n1653), .QN(
        n5069) );
  OAI22X1 U6089 ( .IN1(n6182), .IN2(n5715), .IN3(n5725), .IN4(n1648), .QN(
        n5070) );
  OAI22X1 U6090 ( .IN1(n6181), .IN2(n5715), .IN3(n5724), .IN4(n1643), .QN(
        n5071) );
  OAI22X1 U6091 ( .IN1(n6180), .IN2(n5715), .IN3(n5724), .IN4(n1638), .QN(
        n5072) );
  OAI22X1 U6092 ( .IN1(n6179), .IN2(n5715), .IN3(n5724), .IN4(n1633), .QN(
        n5073) );
  OAI22X1 U6093 ( .IN1(n6178), .IN2(n5715), .IN3(n5724), .IN4(n1628), .QN(
        n5074) );
  OAI22X1 U6094 ( .IN1(n6177), .IN2(n5715), .IN3(n5724), .IN4(n1623), .QN(
        n5075) );
  OAI22X1 U6095 ( .IN1(n6176), .IN2(n5714), .IN3(n5723), .IN4(n1618), .QN(
        n5076) );
  OAI22X1 U6096 ( .IN1(n6175), .IN2(n5714), .IN3(n5723), .IN4(n1613), .QN(
        n5077) );
  OAI22X1 U6097 ( .IN1(n6174), .IN2(n5714), .IN3(n5723), .IN4(n1608), .QN(
        n5078) );
  OAI22X1 U6098 ( .IN1(n6173), .IN2(n5712), .IN3(n5723), .IN4(n1603), .QN(
        n5079) );
  OAI22X1 U6099 ( .IN1(n6172), .IN2(n5714), .IN3(n5723), .IN4(n1598), .QN(
        n5080) );
  OAI22X1 U6100 ( .IN1(n6171), .IN2(n5714), .IN3(n5719), .IN4(n1593), .QN(
        n5081) );
  OAI22X1 U6101 ( .IN1(n6170), .IN2(n5714), .IN3(n5719), .IN4(n1588), .QN(
        n5082) );
  OAI22X1 U6102 ( .IN1(n6169), .IN2(n5714), .IN3(n5723), .IN4(n1583), .QN(
        n5083) );
  OAI22X1 U6103 ( .IN1(n6168), .IN2(n5714), .IN3(n4910), .IN4(n1578), .QN(
        n5084) );
  OAI22X1 U6104 ( .IN1(n6167), .IN2(n5714), .IN3(n5725), .IN4(n1573), .QN(
        n5085) );
  OAI22X1 U6105 ( .IN1(n6166), .IN2(n5714), .IN3(n5722), .IN4(n1568), .QN(
        n5086) );
  OAI22X1 U6106 ( .IN1(n5708), .IN2(n6217), .IN3(n5720), .IN4(n1163), .QN(
        n5087) );
  OAI22X1 U6107 ( .IN1(n5710), .IN2(n5855), .IN3(n5721), .IN4(n1143), .QN(
        n5088) );
  OAI22X1 U6108 ( .IN1(n5286), .IN2(n4093), .IN3(n5855), .IN4(n5299), .QN(
        n5089) );
  OAI22X1 U6109 ( .IN1(n5286), .IN2(n4109), .IN3(n6217), .IN4(n5297), .QN(
        n5090) );
  OAI22X1 U6110 ( .IN1(n5295), .IN2(n4557), .IN3(n6165), .IN4(n5303), .QN(
        n5091) );
  OAI22X1 U6111 ( .IN1(n5295), .IN2(n4553), .IN3(n6164), .IN4(n5303), .QN(
        n5092) );
  OAI22X1 U6112 ( .IN1(n5295), .IN2(n4549), .IN3(n6163), .IN4(n5303), .QN(
        n5093) );
  OAI22X1 U6113 ( .IN1(n5295), .IN2(n4545), .IN3(n6162), .IN4(n5303), .QN(
        n5094) );
  OAI22X1 U6114 ( .IN1(n5295), .IN2(n4541), .IN3(n6161), .IN4(n5303), .QN(
        n5095) );
  OAI22X1 U6115 ( .IN1(n5295), .IN2(n4537), .IN3(n6192), .IN4(n5303), .QN(
        n5096) );
  OAI22X1 U6116 ( .IN1(n5295), .IN2(n4533), .IN3(n6191), .IN4(n5303), .QN(
        n5097) );
  OAI22X1 U6117 ( .IN1(n5295), .IN2(n4529), .IN3(n6190), .IN4(n5303), .QN(
        n5098) );
  OAI22X1 U6118 ( .IN1(n5295), .IN2(n4525), .IN3(n6189), .IN4(n5303), .QN(
        n5099) );
  OAI22X1 U6119 ( .IN1(n5294), .IN2(n4521), .IN3(n6188), .IN4(n5303), .QN(
        n5100) );
  OAI22X1 U6120 ( .IN1(n5294), .IN2(n4517), .IN3(n6187), .IN4(n5302), .QN(
        n5101) );
  OAI22X1 U6121 ( .IN1(n5294), .IN2(n4513), .IN3(n6186), .IN4(n5302), .QN(
        n5102) );
  OAI22X1 U6122 ( .IN1(n5294), .IN2(n4509), .IN3(n6185), .IN4(n5302), .QN(
        n5103) );
  OAI22X1 U6123 ( .IN1(n5294), .IN2(n4505), .IN3(n6184), .IN4(n5302), .QN(
        n5104) );
  OAI22X1 U6124 ( .IN1(n5294), .IN2(n4501), .IN3(n6183), .IN4(n5302), .QN(
        n5105) );
  OAI22X1 U6125 ( .IN1(n5294), .IN2(n4497), .IN3(n6182), .IN4(n5302), .QN(
        n5106) );
  OAI22X1 U6126 ( .IN1(n5294), .IN2(n4493), .IN3(n6181), .IN4(n5302), .QN(
        n5107) );
  OAI22X1 U6127 ( .IN1(n5294), .IN2(n4489), .IN3(n6180), .IN4(n5302), .QN(
        n5108) );
  OAI22X1 U6128 ( .IN1(n5294), .IN2(n4485), .IN3(n6179), .IN4(n5302), .QN(
        n5109) );
  OAI22X1 U6129 ( .IN1(n5294), .IN2(n4481), .IN3(n6178), .IN4(n5302), .QN(
        n5110) );
  OAI22X1 U6130 ( .IN1(n5294), .IN2(n4477), .IN3(n6177), .IN4(n5302), .QN(
        n5111) );
  OAI22X1 U6131 ( .IN1(n5293), .IN2(n4473), .IN3(n6176), .IN4(n5302), .QN(
        n5112) );
  OAI22X1 U6132 ( .IN1(n5293), .IN2(n4469), .IN3(n6175), .IN4(n5302), .QN(
        n5113) );
  OAI22X1 U6133 ( .IN1(n5293), .IN2(n4465), .IN3(n6174), .IN4(n5302), .QN(
        n5114) );
  OAI22X1 U6134 ( .IN1(n5293), .IN2(n4461), .IN3(n6173), .IN4(n5302), .QN(
        n5115) );
  OAI22X1 U6135 ( .IN1(n5293), .IN2(n4457), .IN3(n6172), .IN4(n5301), .QN(
        n5116) );
  OAI22X1 U6136 ( .IN1(n5293), .IN2(n4453), .IN3(n6171), .IN4(n5301), .QN(
        n5117) );
  OAI22X1 U6137 ( .IN1(n5293), .IN2(n4449), .IN3(n6170), .IN4(n5301), .QN(
        n5118) );
  OAI22X1 U6138 ( .IN1(n5293), .IN2(n4445), .IN3(n6169), .IN4(n5301), .QN(
        n5119) );
  OAI22X1 U6139 ( .IN1(n5293), .IN2(n4441), .IN3(n6168), .IN4(n5301), .QN(
        n5120) );
  OAI22X1 U6140 ( .IN1(n5293), .IN2(n4437), .IN3(n6167), .IN4(n5301), .QN(
        n5121) );
  OAI22X1 U6141 ( .IN1(n5293), .IN2(n4433), .IN3(n6166), .IN4(n5301), .QN(
        n5122) );
  OAI22X1 U6142 ( .IN1(n5795), .IN2(n4598), .IN3(n5801), .IN4(n5855), .QN(
        n5123) );
  OAI22X1 U6143 ( .IN1(n5796), .IN2(n4614), .IN3(n5802), .IN4(n6217), .QN(
        n5124) );
  OAI22X1 U6144 ( .IN1(n5795), .IN2(n1093), .IN3(n5800), .IN4(n6165), .QN(
        n5125) );
  OAI22X1 U6145 ( .IN1(n5795), .IN2(n1089), .IN3(n5800), .IN4(n6164), .QN(
        n5126) );
  OAI22X1 U6146 ( .IN1(n5795), .IN2(n1085), .IN3(n5800), .IN4(n6163), .QN(
        n5127) );
  OAI22X1 U6147 ( .IN1(n5795), .IN2(n1081), .IN3(n5806), .IN4(n6162), .QN(
        n5128) );
  OAI22X1 U6148 ( .IN1(n5795), .IN2(n1077), .IN3(n5789), .IN4(n6161), .QN(
        n5129) );
  OAI22X1 U6149 ( .IN1(n5795), .IN2(n1073), .IN3(n5788), .IN4(n6192), .QN(
        n5130) );
  OAI22X1 U6150 ( .IN1(n5794), .IN2(n1069), .IN3(n5787), .IN4(n6191), .QN(
        n5131) );
  OAI22X1 U6151 ( .IN1(n5794), .IN2(n1065), .IN3(n5805), .IN4(n6190), .QN(
        n5132) );
  OAI22X1 U6152 ( .IN1(n5794), .IN2(n1061), .IN3(n5800), .IN4(n6189), .QN(
        n5133) );
  OAI22X1 U6153 ( .IN1(n5794), .IN2(n1057), .IN3(n5805), .IN4(n6188), .QN(
        n5134) );
  OAI22X1 U6154 ( .IN1(n5794), .IN2(n1053), .IN3(n5804), .IN4(n6187), .QN(
        n5135) );
  OAI22X1 U6155 ( .IN1(n5794), .IN2(n1049), .IN3(n5803), .IN4(n6186), .QN(
        n5136) );
  OAI22X1 U6156 ( .IN1(n5794), .IN2(n1045), .IN3(n5804), .IN4(n6185), .QN(
        n5137) );
  OAI22X1 U6157 ( .IN1(n5794), .IN2(n1041), .IN3(n5800), .IN4(n6184), .QN(
        n5138) );
  OAI22X1 U6158 ( .IN1(n5794), .IN2(n1037), .IN3(n5807), .IN4(n6183), .QN(
        n5139) );
  OAI22X1 U6159 ( .IN1(n5794), .IN2(n1033), .IN3(n5805), .IN4(n6182), .QN(
        n5140) );
  OAI22X1 U6160 ( .IN1(n5794), .IN2(n1029), .IN3(n5804), .IN4(n6181), .QN(
        n5141) );
  OAI22X1 U6161 ( .IN1(n5794), .IN2(n1025), .IN3(n5802), .IN4(n6180), .QN(
        n5142) );
  OAI22X1 U6162 ( .IN1(n5793), .IN2(n1021), .IN3(n5801), .IN4(n6179), .QN(
        n5143) );
  OAI22X1 U6163 ( .IN1(n5793), .IN2(n1017), .IN3(n5806), .IN4(n6178), .QN(
        n5144) );
  OAI22X1 U6164 ( .IN1(n5793), .IN2(n1013), .IN3(n5805), .IN4(n6177), .QN(
        n5145) );
  OAI22X1 U6165 ( .IN1(n5793), .IN2(n1009), .IN3(n5801), .IN4(n6176), .QN(
        n5146) );
  OAI22X1 U6166 ( .IN1(n5793), .IN2(n1005), .IN3(n5807), .IN4(n6175), .QN(
        n5147) );
  OAI22X1 U6167 ( .IN1(n5793), .IN2(n1001), .IN3(n5804), .IN4(n6174), .QN(
        n5148) );
  OAI22X1 U6168 ( .IN1(n5793), .IN2(n997), .IN3(n5806), .IN4(n6173), .QN(n5149) );
  OAI22X1 U6169 ( .IN1(n5793), .IN2(n993), .IN3(n5802), .IN4(n6172), .QN(n5150) );
  OAI22X1 U6170 ( .IN1(n5793), .IN2(n989), .IN3(n5803), .IN4(n6171), .QN(n5151) );
  OAI22X1 U6171 ( .IN1(n5793), .IN2(n985), .IN3(n5804), .IN4(n6170), .QN(n5152) );
  OAI22X1 U6172 ( .IN1(n5793), .IN2(n981), .IN3(n5805), .IN4(n6169), .QN(n5153) );
  OAI22X1 U6173 ( .IN1(n5793), .IN2(n977), .IN3(n5804), .IN4(n6168), .QN(n5154) );
  OAI22X1 U6174 ( .IN1(n5792), .IN2(n973), .IN3(n5803), .IN4(n6167), .QN(n5155) );
  OAI22X1 U6175 ( .IN1(n5792), .IN2(n969), .IN3(n5807), .IN4(n6166), .QN(n5156) );
  OAI22X1 U6176 ( .IN1(n6165), .IN2(n5716), .IN3(n5726), .IN4(n1723), .QN(
        n5157) );
  OAI22X1 U6177 ( .IN1(n6164), .IN2(n5716), .IN3(n5722), .IN4(n1718), .QN(
        n5158) );
  OAI22X1 U6178 ( .IN1(n6163), .IN2(n5716), .IN3(n5721), .IN4(n1713), .QN(
        n5159) );
  OAI22X1 U6179 ( .IN1(n6162), .IN2(n5716), .IN3(n5719), .IN4(n1708), .QN(
        n5160) );
  OAI22X1 U6180 ( .IN1(n6161), .IN2(n5716), .IN3(n5720), .IN4(n1703), .QN(
        n5161) );
  OAI22X1 U6181 ( .IN1(n6192), .IN2(n5716), .IN3(n5718), .IN4(n1698), .QN(
        n5162) );
  OAI22X1 U6182 ( .IN1(n6191), .IN2(n5716), .IN3(n5726), .IN4(n1693), .QN(
        n5163) );
  AND2X1 U6183 ( .IN1(\decodedPacket[4][5] ), .IN2(n5268), .Q(n5164) );
  AND2X1 U6184 ( .IN1(\decodedPacket[4][6] ), .IN2(n5268), .Q(n5165) );
  AND2X1 U6185 ( .IN1(\decodedPacket[4][7] ), .IN2(n5268), .Q(n5166) );
  AND2X1 U6186 ( .IN1(\decodedPacket[4][8] ), .IN2(n5268), .Q(n5167) );
  AND2X1 U6187 ( .IN1(\decodedPacket[4][9] ), .IN2(n5268), .Q(n5168) );
  AND2X1 U6188 ( .IN1(\decodedPacket[4][10] ), .IN2(n5268), .Q(n5169) );
  AND2X1 U6189 ( .IN1(\decodedPacket[4][12] ), .IN2(n5268), .Q(n5170) );
  AND2X1 U6190 ( .IN1(\decodedPacket[4][5] ), .IN2(n5270), .Q(n5171) );
  AND2X1 U6191 ( .IN1(\decodedPacket[4][6] ), .IN2(n5270), .Q(n5172) );
  AND2X1 U6192 ( .IN1(\decodedPacket[4][7] ), .IN2(n5270), .Q(n5173) );
  AND2X1 U6193 ( .IN1(\decodedPacket[4][8] ), .IN2(n5270), .Q(n5174) );
  AND2X1 U6194 ( .IN1(\decodedPacket[4][9] ), .IN2(n5270), .Q(n5175) );
  AND2X1 U6195 ( .IN1(\decodedPacket[4][10] ), .IN2(n5270), .Q(n5176) );
  AND2X1 U6196 ( .IN1(\decodedPacket[4][12] ), .IN2(n5270), .Q(n5177) );
  AND2X1 U6197 ( .IN1(\decodedPacket[4][5] ), .IN2(n5272), .Q(n5178) );
  AND2X1 U6198 ( .IN1(\decodedPacket[4][6] ), .IN2(n5272), .Q(n5179) );
  AND2X1 U6199 ( .IN1(\decodedPacket[4][7] ), .IN2(n5272), .Q(n5180) );
  AND2X1 U6200 ( .IN1(\decodedPacket[4][8] ), .IN2(n5272), .Q(n5181) );
  AND2X1 U6201 ( .IN1(\decodedPacket[4][9] ), .IN2(n5272), .Q(n5182) );
  AND2X1 U6202 ( .IN1(\decodedPacket[4][10] ), .IN2(n5272), .Q(n5183) );
  AND2X1 U6203 ( .IN1(\decodedPacket[4][12] ), .IN2(n5272), .Q(n5184) );
  AND2X1 U6204 ( .IN1(\decodedPacket[4][5] ), .IN2(n5274), .Q(n5185) );
  AND2X1 U6205 ( .IN1(\decodedPacket[4][6] ), .IN2(n5274), .Q(n5186) );
  AND2X1 U6206 ( .IN1(\decodedPacket[4][7] ), .IN2(n5274), .Q(n5187) );
  AND2X1 U6207 ( .IN1(\decodedPacket[4][8] ), .IN2(n5274), .Q(n5188) );
  AND2X1 U6208 ( .IN1(\decodedPacket[4][9] ), .IN2(n5274), .Q(n5189) );
  AND2X1 U6209 ( .IN1(\decodedPacket[4][10] ), .IN2(n5274), .Q(n5190) );
  AND2X1 U6210 ( .IN1(\decodedPacket[4][12] ), .IN2(n5274), .Q(n5191) );
  NAND2X1 U6211 ( .IN1(n5696), .IN2(n5195), .QN(n1143) );
  NAND2X1 U6212 ( .IN1(n5616), .IN2(n5196), .QN(n1814) );
  NAND2X1 U6213 ( .IN1(n5616), .IN2(n5197), .QN(n1790) );
  NAND2X1 U6214 ( .IN1(n5696), .IN2(n5198), .QN(n1163) );
  NAND2X1 U6215 ( .IN1(n5617), .IN2(n5202), .QN(n2378) );
  NAND2X1 U6216 ( .IN1(n5617), .IN2(n5203), .QN(n2372) );
  NAND2X1 U6217 ( .IN1(n5617), .IN2(n5204), .QN(n2366) );
  NAND2X1 U6218 ( .IN1(n5617), .IN2(n5205), .QN(n2360) );
  NAND2X1 U6219 ( .IN1(n5616), .IN2(n5206), .QN(n2354) );
  NAND2X1 U6220 ( .IN1(n5616), .IN2(n5207), .QN(n2348) );
  NAND2X1 U6221 ( .IN1(n5616), .IN2(n5208), .QN(n2342) );
  NAND2X1 U6222 ( .IN1(n5616), .IN2(n5209), .QN(n2336) );
  NAND2X1 U6223 ( .IN1(n5616), .IN2(n5210), .QN(n2330) );
  NAND2X1 U6224 ( .IN1(n5616), .IN2(n5211), .QN(n2324) );
  NAND2X1 U6225 ( .IN1(n5616), .IN2(n5212), .QN(n2318) );
  NAND2X1 U6226 ( .IN1(n5616), .IN2(n5213), .QN(n2312) );
  NAND2X1 U6227 ( .IN1(n5616), .IN2(n5214), .QN(n2306) );
  NAND2X1 U6228 ( .IN1(n5616), .IN2(n5215), .QN(n2300) );
  NAND2X1 U6229 ( .IN1(n5618), .IN2(n5216), .QN(n2486) );
  NAND2X1 U6230 ( .IN1(n5618), .IN2(n5217), .QN(n2480) );
  NAND2X1 U6231 ( .IN1(n5618), .IN2(n5218), .QN(n2474) );
  NAND2X1 U6232 ( .IN1(n5618), .IN2(n5219), .QN(n2468) );
  NAND2X1 U6233 ( .IN1(n5618), .IN2(n5220), .QN(n2462) );
  NAND2X1 U6234 ( .IN1(n5618), .IN2(n5221), .QN(n2456) );
  NAND2X1 U6235 ( .IN1(n5618), .IN2(n5222), .QN(n2450) );
  NAND2X1 U6236 ( .IN1(n5618), .IN2(n5223), .QN(n2444) );
  NAND2X1 U6237 ( .IN1(n5618), .IN2(n5224), .QN(n2438) );
  NAND2X1 U6238 ( .IN1(n5618), .IN2(n5225), .QN(n2432) );
  NAND2X1 U6239 ( .IN1(n5617), .IN2(n5226), .QN(n2426) );
  NAND2X1 U6240 ( .IN1(n5617), .IN2(n5227), .QN(n2420) );
  NAND2X1 U6241 ( .IN1(n5617), .IN2(n5228), .QN(n2414) );
  NAND2X1 U6242 ( .IN1(n5617), .IN2(n5229), .QN(n2408) );
  NAND2X1 U6243 ( .IN1(n5617), .IN2(n5230), .QN(n2402) );
  NAND2X1 U6244 ( .IN1(n5617), .IN2(n5231), .QN(n2396) );
  NAND2X1 U6245 ( .IN1(n5617), .IN2(n5232), .QN(n2390) );
  NAND2X1 U6246 ( .IN1(n5617), .IN2(n5233), .QN(n2384) );
  NAND2X1 U6247 ( .IN1(n5698), .IN2(n5234), .QN(n1688) );
  NAND2X1 U6248 ( .IN1(n5698), .IN2(n5235), .QN(n1683) );
  NAND2X1 U6249 ( .IN1(n5698), .IN2(n5236), .QN(n1678) );
  NAND2X1 U6250 ( .IN1(n5697), .IN2(n5237), .QN(n1673) );
  NAND2X1 U6251 ( .IN1(n5697), .IN2(n5238), .QN(n1668) );
  NAND2X1 U6252 ( .IN1(n5697), .IN2(n5239), .QN(n1663) );
  NAND2X1 U6253 ( .IN1(n5697), .IN2(n5240), .QN(n1658) );
  NAND2X1 U6254 ( .IN1(n5697), .IN2(n5241), .QN(n1653) );
  NAND2X1 U6255 ( .IN1(n5697), .IN2(n5242), .QN(n1648) );
  NAND2X1 U6256 ( .IN1(n5697), .IN2(n5243), .QN(n1643) );
  NAND2X1 U6257 ( .IN1(n5697), .IN2(n5244), .QN(n1638) );
  NAND2X1 U6258 ( .IN1(n5697), .IN2(n5245), .QN(n1633) );
  NAND2X1 U6259 ( .IN1(n5697), .IN2(n5246), .QN(n1628) );
  NAND2X1 U6260 ( .IN1(n5697), .IN2(n5247), .QN(n1623) );
  NAND2X1 U6261 ( .IN1(n5697), .IN2(n5248), .QN(n1618) );
  NAND2X1 U6262 ( .IN1(n5696), .IN2(n5249), .QN(n1613) );
  NAND2X1 U6263 ( .IN1(n5696), .IN2(n5250), .QN(n1608) );
  NAND2X1 U6264 ( .IN1(n5696), .IN2(n5251), .QN(n1603) );
  NAND2X1 U6265 ( .IN1(n5696), .IN2(n5252), .QN(n1598) );
  NAND2X1 U6266 ( .IN1(n5696), .IN2(n5253), .QN(n1593) );
  NAND2X1 U6267 ( .IN1(n5696), .IN2(n5254), .QN(n1588) );
  NAND2X1 U6268 ( .IN1(n5696), .IN2(n5255), .QN(n1583) );
  NAND2X1 U6269 ( .IN1(n5696), .IN2(n5256), .QN(n1578) );
  NAND2X1 U6270 ( .IN1(n5696), .IN2(n5257), .QN(n1573) );
  NAND2X1 U6271 ( .IN1(n5696), .IN2(n5258), .QN(n1568) );
  NAND2X1 U6272 ( .IN1(n5698), .IN2(n5259), .QN(n1723) );
  NAND2X1 U6273 ( .IN1(n5698), .IN2(n5260), .QN(n1718) );
  NAND2X1 U6274 ( .IN1(n5698), .IN2(n5261), .QN(n1713) );
  NAND2X1 U6275 ( .IN1(n5698), .IN2(n5262), .QN(n1708) );
  NAND2X1 U6276 ( .IN1(n5698), .IN2(n5263), .QN(n1703) );
  NAND2X1 U6277 ( .IN1(n5698), .IN2(n5264), .QN(n1698) );
  NAND2X1 U6278 ( .IN1(n5698), .IN2(n5265), .QN(n1693) );
  NAND2X1 U6279 ( .IN1(N6449), .IN2(\add_177_I7_aco/carry[5] ), .QN(n5192) );
  OR2X1 U6280 ( .IN1(N4311), .IN2(N4312), .Q(n5193) );
  OR3X1 U6281 ( .IN1(N6447), .IN2(N6449), .IN3(N6448), .Q(n5194) );
  INVX0 U6282 ( .INP(\decodedPacket[3][74] ), .ZN(n6088) );
  INVX0 U6283 ( .INP(\decodedPacket[3][76] ), .ZN(n6089) );
  INVX0 U6284 ( .INP(\decodedPacket[3][77] ), .ZN(n6090) );
  INVX0 U6285 ( .INP(\decodedPacket[5][74] ), .ZN(n6241) );
  INVX0 U6286 ( .INP(\decodedPacket[5][76] ), .ZN(n6243) );
  INVX0 U6287 ( .INP(\decodedPacket[5][77] ), .ZN(n6244) );
  INVX0 U6288 ( .INP(\decodedPacket[3][73] ), .ZN(n6087) );
  INVX0 U6289 ( .INP(\decodedPacket[3][115] ), .ZN(n6091) );
  INVX0 U6290 ( .INP(\decodedPacket[5][75] ), .ZN(n6242) );
  INVX0 U6291 ( .INP(\decodedPacket[5][115] ), .ZN(n6245) );
  INVX0 U6292 ( .INP(\decodedPacket[7][76] ), .ZN(n6398) );
  INVX0 U6293 ( .INP(\decodedPacket[7][74] ), .ZN(n6396) );
  INVX0 U6294 ( .INP(\decodedPacket[7][77] ), .ZN(n6399) );
  INVX0 U6295 ( .INP(\decodedPacket[7][69] ), .ZN(n6395) );
  INVX0 U6296 ( .INP(\decodedPacket[7][75] ), .ZN(n6397) );
  NBUFFX2 U6297 ( .INP(n5352), .Z(n5268) );
  NBUFFX2 U6298 ( .INP(n5411), .Z(n5270) );
  NBUFFX2 U6299 ( .INP(n5470), .Z(n5272) );
  NBUFFX2 U6300 ( .INP(n5529), .Z(n5274) );
  NBUFFX2 U6301 ( .INP(n5352), .Z(n5269) );
  NBUFFX2 U6302 ( .INP(n5411), .Z(n5271) );
  NBUFFX2 U6303 ( .INP(n5470), .Z(n5273) );
  NBUFFX2 U6304 ( .INP(n5529), .Z(n5275) );
  NOR2X0 U6305 ( .IN1(n4066), .IN2(N8582), .QN(n1752) );
  NOR2X0 U6306 ( .IN1(n5982), .IN2(n4066), .QN(n2909) );
  INVX0 U6307 ( .INP(N8582), .ZN(n5982) );
  NOR2X0 U6308 ( .IN1(N2175), .IN2(N2174), .QN(n1754) );
  NOR2X0 U6309 ( .IN1(n5984), .IN2(n5193), .QN(n2907) );
  INVX0 U6310 ( .INP(N4310), .ZN(n5984) );
  NOR2X0 U6311 ( .IN1(n5193), .IN2(N4310), .QN(n1755) );
  NOR2X0 U6312 ( .IN1(n5194), .IN2(N6446), .QN(n1753) );
  NOR2X0 U6313 ( .IN1(n5983), .IN2(n5194), .QN(n2910) );
  INVX0 U6314 ( .INP(N6446), .ZN(n5983) );
  NOR2X0 U6315 ( .IN1(n5985), .IN2(N2175), .QN(n2908) );
  INVX0 U6316 ( .INP(N2174), .ZN(n5985) );
  NOR2X0 U6317 ( .IN1(n1140), .IN2(n5761), .QN(N9922) );
  NAND2X1 U6318 ( .IN1(n5727), .IN2(n5088), .QN(n1141) );
  NOR2X0 U6319 ( .IN1(n3696), .IN2(n5399), .QN(N10312) );
  NAND2X1 U6320 ( .IN1(n5363), .IN2(n4988), .QN(n3697) );
  NOR2X0 U6321 ( .IN1(n3312), .IN2(n5458), .QN(N10442) );
  NAND2X1 U6322 ( .IN1(n5422), .IN2(n4989), .QN(n3313) );
  NOR2X0 U6323 ( .IN1(n2928), .IN2(n5517), .QN(N10572) );
  NAND2X1 U6324 ( .IN1(n5481), .IN2(n4990), .QN(n2929) );
  NOR2X0 U6325 ( .IN1(n2539), .IN2(n5576), .QN(N10702) );
  NAND2X1 U6326 ( .IN1(n5539), .IN2(n4991), .QN(n2540) );
  NOR2X0 U6327 ( .IN1(n1787), .IN2(n5671), .QN(N9792) );
  NAND2X1 U6328 ( .IN1(n5637), .IN2(n5042), .QN(n1788) );
  NOR2X0 U6329 ( .IN1(n4090), .IN2(n5338), .QN(N10182) );
  NAND2X1 U6330 ( .IN1(n5304), .IN2(n5089), .QN(n4091) );
  NOR2X0 U6331 ( .IN1(n4595), .IN2(n5843), .QN(N10052) );
  NAND2X1 U6332 ( .IN1(n5808), .IN2(n5123), .QN(n4596) );
  NAND2X1 U6333 ( .IN1(\decodedPacket[0][121] ), .IN2(n5586), .QN(n1792) );
  INVX0 U6334 ( .INP(\decodedPacket[3][119] ), .ZN(n6068) );
  INVX0 U6335 ( .INP(\decodedPacket[5][119] ), .ZN(n6222) );
  NBUFFX2 U6336 ( .INP(decodedVector_o[3]), .Z(n5887) );
  NBUFFX2 U6337 ( .INP(decodedVector_o[3]), .Z(n5888) );
  NBUFFX2 U6338 ( .INP(decodedVector_o[3]), .Z(n5889) );
  NBUFFX2 U6339 ( .INP(decodedVector_o[3]), .Z(n5890) );
  NBUFFX2 U6340 ( .INP(decodedVector_o[3]), .Z(n5891) );
  NBUFFX2 U6341 ( .INP(decodedVector_o[3]), .Z(n5892) );
  NBUFFX2 U6342 ( .INP(decodedVector_o[3]), .Z(n5893) );
  NBUFFX2 U6343 ( .INP(decodedVector_o[3]), .Z(n5894) );
  NBUFFX2 U6344 ( .INP(decodedVector_o[3]), .Z(n5895) );
  NBUFFX2 U6345 ( .INP(decodedVector_o[3]), .Z(n5896) );
  NBUFFX2 U6346 ( .INP(decodedVector_o[1]), .Z(n5867) );
  NBUFFX2 U6347 ( .INP(decodedVector_o[1]), .Z(n5868) );
  NBUFFX2 U6348 ( .INP(decodedVector_o[1]), .Z(n5869) );
  NBUFFX2 U6349 ( .INP(decodedVector_o[1]), .Z(n5870) );
  NBUFFX2 U6350 ( .INP(decodedVector_o[1]), .Z(n5871) );
  NBUFFX2 U6351 ( .INP(decodedVector_o[1]), .Z(n5872) );
  NBUFFX2 U6352 ( .INP(decodedVector_o[1]), .Z(n5873) );
  NBUFFX2 U6353 ( .INP(decodedVector_o[1]), .Z(n5874) );
  NBUFFX2 U6354 ( .INP(decodedVector_o[1]), .Z(n5875) );
  NBUFFX2 U6355 ( .INP(decodedVector_o[1]), .Z(n5876) );
  INVX0 U6356 ( .INP(\decodedPacket[7][119] ), .ZN(n6376) );
  INVX0 U6357 ( .INP(\decodedPacket[3][70] ), .ZN(n6042) );
  INVX0 U6358 ( .INP(\decodedPacket[5][70] ), .ZN(n6196) );
  INVX0 U6359 ( .INP(\decodedPacket[3][91] ), .ZN(n6075) );
  INVX0 U6360 ( .INP(\decodedPacket[5][91] ), .ZN(n6229) );
  INVX0 U6361 ( .INP(\decodedPacket[3][116] ), .ZN(n6065) );
  INVX0 U6362 ( .INP(\decodedPacket[5][116] ), .ZN(n6219) );
  INVX0 U6363 ( .INP(\decodedPacket[3][98] ), .ZN(n6064) );
  INVX0 U6364 ( .INP(\decodedPacket[7][70] ), .ZN(n6350) );
  INVX0 U6365 ( .INP(\decodedPacket[5][98] ), .ZN(n6218) );
  INVX0 U6366 ( .INP(\decodedPacket[7][116] ), .ZN(n6373) );
  INVX0 U6367 ( .INP(\decodedPacket[7][91] ), .ZN(n6383) );
  INVX0 U6368 ( .INP(\decodedPacket[7][98] ), .ZN(n6372) );
  AND2X1 U6369 ( .IN1(\decodedPacket[2][121] ), .IN2(n5691), .Q(n5195) );
  INVX0 U6370 ( .INP(\decodedPacket[4][121] ), .ZN(n5855) );
  NAND2X1 U6371 ( .IN1(n5773), .IN2(\decodedPacket[2][121] ), .QN(n4598) );
  NAND2X1 U6372 ( .IN1(n5276), .IN2(\decodedPacket[2][121] ), .QN(n4093) );
  INVX0 U6373 ( .INP(\decodedPacket[2][84] ), .ZN(n6045) );
  INVX0 U6374 ( .INP(\decodedPacket[2][77] ), .ZN(n6044) );
  INVX0 U6375 ( .INP(\decodedPacket[2][119] ), .ZN(n6040) );
  NOR2X0 U6376 ( .IN1(n5340), .IN2(n5282), .QN(n4578) );
  INVX0 U6377 ( .INP(N2173), .ZN(n5990) );
  NOR4X0 U6378 ( .IN1(\add_177_I3_aco/A[1] ), .IN2(n5763), .IN3(n5693), .IN4(
        n5702), .QN(n1750) );
  INVX0 U6379 ( .INP(N1069), .ZN(n5991) );
  INVX0 U6380 ( .INP(N1070), .ZN(n5986) );
  INVX0 U6381 ( .INP(N8581), .ZN(n5987) );
  INVX0 U6382 ( .INP(N4309), .ZN(n5989) );
  INVX0 U6383 ( .INP(N6445), .ZN(n5988) );
  NOR2X0 U6384 ( .IN1(n1160), .IN2(n5761), .QN(N9918) );
  NAND2X1 U6385 ( .IN1(n5727), .IN2(n5087), .QN(n1161) );
  NOR2X0 U6386 ( .IN1(n3708), .IN2(n5399), .QN(N10308) );
  NAND2X1 U6387 ( .IN1(n5363), .IN2(n4992), .QN(n3709) );
  NOR2X0 U6388 ( .IN1(n3324), .IN2(n5458), .QN(N10438) );
  NAND2X1 U6389 ( .IN1(n5422), .IN2(n4993), .QN(n3325) );
  NOR2X0 U6390 ( .IN1(n2940), .IN2(n5517), .QN(N10568) );
  NAND2X1 U6391 ( .IN1(n5481), .IN2(n4994), .QN(n2941) );
  NOR2X0 U6392 ( .IN1(n2551), .IN2(n5576), .QN(N10698) );
  NAND2X1 U6393 ( .IN1(n5539), .IN2(n4933), .QN(n2552) );
  NOR2X0 U6394 ( .IN1(n1811), .IN2(n5671), .QN(N9788) );
  NAND2X1 U6395 ( .IN1(n5637), .IN2(n5043), .QN(n1812) );
  NOR2X0 U6396 ( .IN1(n4106), .IN2(n5338), .QN(N10178) );
  NAND2X1 U6397 ( .IN1(n5304), .IN2(n5090), .QN(n4107) );
  NOR2X0 U6398 ( .IN1(n4611), .IN2(n5843), .QN(N10048) );
  NAND2X1 U6399 ( .IN1(n5808), .IN2(n5124), .QN(n4612) );
  INVX0 U6400 ( .INP(\decodedPacket[3][120] ), .ZN(n6076) );
  INVX0 U6401 ( .INP(\decodedPacket[5][120] ), .ZN(n6230) );
  INVX0 U6402 ( .INP(\decodedPacket[4][98] ), .ZN(n6152) );
  INVX0 U6403 ( .INP(\decodedPacket[6][98] ), .ZN(n6306) );
  INVX0 U6404 ( .INP(\decodedPacket[4][84] ), .ZN(n6199) );
  INVX0 U6405 ( .INP(\decodedPacket[6][84] ), .ZN(n6353) );
  INVX0 U6406 ( .INP(\decodedPacket[7][120] ), .ZN(n6384) );
  INVX0 U6407 ( .INP(\decodedPacket[4][77] ), .ZN(n6198) );
  INVX0 U6408 ( .INP(\decodedPacket[6][77] ), .ZN(n6352) );
  INVX0 U6409 ( .INP(\decodedPacket[4][119] ), .ZN(n6194) );
  INVX0 U6410 ( .INP(\decodedPacket[6][119] ), .ZN(n6348) );
  NBUFFX2 U6411 ( .INP(n5407), .Z(n5404) );
  NBUFFX2 U6412 ( .INP(n5404), .Z(n5405) );
  NBUFFX2 U6413 ( .INP(n5409), .Z(n5406) );
  NBUFFX2 U6414 ( .INP(n5397), .Z(n5407) );
  NBUFFX2 U6415 ( .INP(n5457), .Z(n5463) );
  NBUFFX2 U6416 ( .INP(n5456), .Z(n5464) );
  NBUFFX2 U6417 ( .INP(n5456), .Z(n5465) );
  NBUFFX2 U6418 ( .INP(n5456), .Z(n5466) );
  NBUFFX2 U6419 ( .INP(n5515), .Z(n5522) );
  NBUFFX2 U6420 ( .INP(n5515), .Z(n5523) );
  NBUFFX2 U6421 ( .INP(n5515), .Z(n5524) );
  NBUFFX2 U6422 ( .INP(n5515), .Z(n5525) );
  NBUFFX2 U6423 ( .INP(n5573), .Z(n5581) );
  NBUFFX2 U6424 ( .INP(n5574), .Z(n5582) );
  NBUFFX2 U6425 ( .INP(n5574), .Z(n5583) );
  NBUFFX2 U6426 ( .INP(n5398), .Z(n5408) );
  NBUFFX2 U6427 ( .INP(n5457), .Z(n5467) );
  NBUFFX2 U6428 ( .INP(n5516), .Z(n5526) );
  NBUFFX2 U6429 ( .INP(n5575), .Z(n5584) );
  NBUFFX2 U6430 ( .INP(n1757), .Z(n5676) );
  NBUFFX2 U6431 ( .INP(n5679), .Z(n5677) );
  NBUFFX2 U6432 ( .INP(n1757), .Z(n5678) );
  NBUFFX2 U6433 ( .INP(n5676), .Z(n5679) );
  NBUFFX2 U6434 ( .INP(n5679), .Z(n5680) );
  NBUFFX2 U6435 ( .INP(n5678), .Z(n5681) );
  NBUFFX2 U6436 ( .INP(n1757), .Z(n5682) );
  NBUFFX2 U6437 ( .INP(n4070), .Z(n5343) );
  NBUFFX2 U6438 ( .INP(n4070), .Z(n5344) );
  NBUFFX2 U6439 ( .INP(n4070), .Z(n5345) );
  NBUFFX2 U6440 ( .INP(n4070), .Z(n5346) );
  NBUFFX2 U6441 ( .INP(n4070), .Z(n5347) );
  NBUFFX2 U6442 ( .INP(n4070), .Z(n5348) );
  NBUFFX2 U6443 ( .INP(n4070), .Z(n5349) );
  NBUFFX2 U6444 ( .INP(n4070), .Z(n5350) );
  NBUFFX2 U6445 ( .INP(n3686), .Z(n5362) );
  NBUFFX2 U6446 ( .INP(n3686), .Z(n5361) );
  NBUFFX2 U6447 ( .INP(n3686), .Z(n5360) );
  NBUFFX2 U6448 ( .INP(n3686), .Z(n5359) );
  NBUFFX2 U6449 ( .INP(n3686), .Z(n5358) );
  NBUFFX2 U6450 ( .INP(n3686), .Z(n5357) );
  NBUFFX2 U6451 ( .INP(n3686), .Z(n5356) );
  NBUFFX2 U6452 ( .INP(n3686), .Z(n5355) );
  NBUFFX2 U6453 ( .INP(n3302), .Z(n5421) );
  NBUFFX2 U6454 ( .INP(n3302), .Z(n5420) );
  NBUFFX2 U6455 ( .INP(n3302), .Z(n5419) );
  NBUFFX2 U6456 ( .INP(n3302), .Z(n5418) );
  NBUFFX2 U6457 ( .INP(n3302), .Z(n5417) );
  NBUFFX2 U6458 ( .INP(n3302), .Z(n5416) );
  NBUFFX2 U6459 ( .INP(n3302), .Z(n5415) );
  NBUFFX2 U6460 ( .INP(n3302), .Z(n5414) );
  NBUFFX2 U6461 ( .INP(n2918), .Z(n5480) );
  NBUFFX2 U6462 ( .INP(n2918), .Z(n5479) );
  NBUFFX2 U6463 ( .INP(n2918), .Z(n5478) );
  NBUFFX2 U6464 ( .INP(n2918), .Z(n5477) );
  NBUFFX2 U6465 ( .INP(n2918), .Z(n5476) );
  NBUFFX2 U6466 ( .INP(n2918), .Z(n5475) );
  NBUFFX2 U6467 ( .INP(n2918), .Z(n5474) );
  NBUFFX2 U6468 ( .INP(n2918), .Z(n5473) );
  NBUFFX2 U6469 ( .INP(n2529), .Z(n5538) );
  NBUFFX2 U6470 ( .INP(n2529), .Z(n5537) );
  NBUFFX2 U6471 ( .INP(n2529), .Z(n5536) );
  NBUFFX2 U6472 ( .INP(n2529), .Z(n5535) );
  NBUFFX2 U6473 ( .INP(n2529), .Z(n5534) );
  NBUFFX2 U6474 ( .INP(n2529), .Z(n5533) );
  NBUFFX2 U6475 ( .INP(n2529), .Z(n5532) );
  NBUFFX2 U6476 ( .INP(n1124), .Z(n5683) );
  NBUFFX2 U6477 ( .INP(n1124), .Z(n5684) );
  NBUFFX2 U6478 ( .INP(n1124), .Z(n5685) );
  NBUFFX2 U6479 ( .INP(n1124), .Z(n5686) );
  NBUFFX2 U6480 ( .INP(n1124), .Z(n5687) );
  NBUFFX2 U6481 ( .INP(n1124), .Z(n5688) );
  NBUFFX2 U6482 ( .INP(n1124), .Z(n5689) );
  NBUFFX2 U6483 ( .INP(n5615), .Z(n5608) );
  NBUFFX2 U6484 ( .INP(n5597), .Z(n5609) );
  NBUFFX2 U6485 ( .INP(n5597), .Z(n5610) );
  NBUFFX2 U6486 ( .INP(n5597), .Z(n5611) );
  NBUFFX2 U6487 ( .INP(n5598), .Z(n5612) );
  NBUFFX2 U6488 ( .INP(n5599), .Z(n5613) );
  NBUFFX2 U6489 ( .INP(n5599), .Z(n5614) );
  NBUFFX2 U6490 ( .INP(n5599), .Z(n5615) );
  NBUFFX2 U6491 ( .INP(n5398), .Z(n5409) );
  NBUFFX2 U6492 ( .INP(n5457), .Z(n5468) );
  NBUFFX2 U6493 ( .INP(n5516), .Z(n5527) );
  NBUFFX2 U6494 ( .INP(n5575), .Z(n5585) );
  NBUFFX2 U6495 ( .INP(n5781), .Z(n5782) );
  NBUFFX2 U6496 ( .INP(n5780), .Z(n5786) );
  NBUFFX2 U6497 ( .INP(n5779), .Z(n5785) );
  NBUFFX2 U6498 ( .INP(n5780), .Z(n5784) );
  NBUFFX2 U6499 ( .INP(n5779), .Z(n5783) );
  NBUFFX2 U6500 ( .INP(n5645), .Z(n5650) );
  NBUFFX2 U6501 ( .INP(n5644), .Z(n5649) );
  NBUFFX2 U6502 ( .INP(n5643), .Z(n5648) );
  NBUFFX2 U6503 ( .INP(n5649), .Z(n5647) );
  NBUFFX2 U6504 ( .INP(n5645), .Z(n5646) );
  NBUFFX2 U6505 ( .INP(n5815), .Z(n5816) );
  NBUFFX2 U6506 ( .INP(n5820), .Z(n5821) );
  NBUFFX2 U6507 ( .INP(n5814), .Z(n5820) );
  NBUFFX2 U6508 ( .INP(n5815), .Z(n5819) );
  NBUFFX2 U6509 ( .INP(n5817), .Z(n5818) );
  NBUFFX2 U6510 ( .INP(n5814), .Z(n5817) );
  NBUFFX2 U6511 ( .INP(n5311), .Z(n5317) );
  NBUFFX2 U6512 ( .INP(n5315), .Z(n5316) );
  NBUFFX2 U6513 ( .INP(n5310), .Z(n5315) );
  NBUFFX2 U6514 ( .INP(n5311), .Z(n5314) );
  NBUFFX2 U6515 ( .INP(n5312), .Z(n5313) );
  NBUFFX2 U6516 ( .INP(n5310), .Z(n5312) );
  NBUFFX2 U6517 ( .INP(n5394), .Z(n5393) );
  NBUFFX2 U6518 ( .INP(n5394), .Z(n5392) );
  NBUFFX2 U6519 ( .INP(n5395), .Z(n5391) );
  NBUFFX2 U6520 ( .INP(n5395), .Z(n5390) );
  NBUFFX2 U6521 ( .INP(n5395), .Z(n5389) );
  NBUFFX2 U6522 ( .INP(n5396), .Z(n5388) );
  NBUFFX2 U6523 ( .INP(n5396), .Z(n5387) );
  NBUFFX2 U6524 ( .INP(n5396), .Z(n5386) );
  NBUFFX2 U6525 ( .INP(n5723), .Z(n5726) );
  NBUFFX2 U6526 ( .INP(n5722), .Z(n5725) );
  NBUFFX2 U6527 ( .INP(n5721), .Z(n5724) );
  NBUFFX2 U6528 ( .INP(n4910), .Z(n5723) );
  NBUFFX2 U6529 ( .INP(n4910), .Z(n5722) );
  NBUFFX2 U6530 ( .INP(n4910), .Z(n5721) );
  NBUFFX2 U6531 ( .INP(n5723), .Z(n5720) );
  NBUFFX2 U6532 ( .INP(n5722), .Z(n5719) );
  NBUFFX2 U6533 ( .INP(n5725), .Z(n5718) );
  NBUFFX2 U6534 ( .INP(n5724), .Z(n5717) );
  NBUFFX2 U6535 ( .INP(n5787), .Z(n5800) );
  NBUFFX2 U6536 ( .INP(n5789), .Z(n5807) );
  NBUFFX2 U6537 ( .INP(n5789), .Z(n5806) );
  NBUFFX2 U6538 ( .INP(n5788), .Z(n5805) );
  NBUFFX2 U6539 ( .INP(n5788), .Z(n5804) );
  NBUFFX2 U6540 ( .INP(n5788), .Z(n5803) );
  NBUFFX2 U6541 ( .INP(n5787), .Z(n5802) );
  NBUFFX2 U6542 ( .INP(n5787), .Z(n5801) );
  NBUFFX2 U6543 ( .INP(n5758), .Z(n5757) );
  NBUFFX2 U6544 ( .INP(n5758), .Z(n5756) );
  NBUFFX2 U6545 ( .INP(n5759), .Z(n5755) );
  NBUFFX2 U6546 ( .INP(n5759), .Z(n5754) );
  NBUFFX2 U6547 ( .INP(n5759), .Z(n5753) );
  NBUFFX2 U6548 ( .INP(n5760), .Z(n5752) );
  NBUFFX2 U6549 ( .INP(n5760), .Z(n5751) );
  NBUFFX2 U6550 ( .INP(n5760), .Z(n5750) );
  NBUFFX2 U6551 ( .INP(n5822), .Z(n5838) );
  NBUFFX2 U6552 ( .INP(n5822), .Z(n5837) );
  NBUFFX2 U6553 ( .INP(n5825), .Z(n5836) );
  NBUFFX2 U6554 ( .INP(n5823), .Z(n5842) );
  NBUFFX2 U6555 ( .INP(n5823), .Z(n5841) );
  NBUFFX2 U6556 ( .INP(n5823), .Z(n5840) );
  NBUFFX2 U6557 ( .INP(n5822), .Z(n5839) );
  NBUFFX2 U6558 ( .INP(n5453), .Z(n5452) );
  NBUFFX2 U6559 ( .INP(n5453), .Z(n5451) );
  NBUFFX2 U6560 ( .INP(n5454), .Z(n5450) );
  NBUFFX2 U6561 ( .INP(n5454), .Z(n5449) );
  NBUFFX2 U6562 ( .INP(n5454), .Z(n5448) );
  NBUFFX2 U6563 ( .INP(n5455), .Z(n5447) );
  NBUFFX2 U6564 ( .INP(n5455), .Z(n5446) );
  NBUFFX2 U6565 ( .INP(n5455), .Z(n5445) );
  NBUFFX2 U6566 ( .INP(n5512), .Z(n5511) );
  NBUFFX2 U6567 ( .INP(n5512), .Z(n5510) );
  NBUFFX2 U6568 ( .INP(n5513), .Z(n5509) );
  NBUFFX2 U6569 ( .INP(n5513), .Z(n5508) );
  NBUFFX2 U6570 ( .INP(n5513), .Z(n5507) );
  NBUFFX2 U6571 ( .INP(n5514), .Z(n5506) );
  NBUFFX2 U6572 ( .INP(n5514), .Z(n5505) );
  NBUFFX2 U6573 ( .INP(n5514), .Z(n5504) );
  NBUFFX2 U6574 ( .INP(n5570), .Z(n5569) );
  NBUFFX2 U6575 ( .INP(n5570), .Z(n5568) );
  NBUFFX2 U6576 ( .INP(n5571), .Z(n5567) );
  NBUFFX2 U6577 ( .INP(n5571), .Z(n5566) );
  NBUFFX2 U6578 ( .INP(n5571), .Z(n5565) );
  NBUFFX2 U6579 ( .INP(n5572), .Z(n5564) );
  NBUFFX2 U6580 ( .INP(n5572), .Z(n5563) );
  NBUFFX2 U6581 ( .INP(n5572), .Z(n5562) );
  NBUFFX2 U6582 ( .INP(n4919), .Z(n5781) );
  NBUFFX2 U6583 ( .INP(n4919), .Z(n5780) );
  NBUFFX2 U6584 ( .INP(n4919), .Z(n5779) );
  NBUFFX2 U6585 ( .INP(n4917), .Z(n5645) );
  NBUFFX2 U6586 ( .INP(n4917), .Z(n5644) );
  NBUFFX2 U6587 ( .INP(n4917), .Z(n5643) );
  NBUFFX2 U6588 ( .INP(n4918), .Z(n5815) );
  NBUFFX2 U6589 ( .INP(n4918), .Z(n5814) );
  NBUFFX2 U6590 ( .INP(n4916), .Z(n5311) );
  NBUFFX2 U6591 ( .INP(n4916), .Z(n5310) );
  INVX0 U6592 ( .INP(\decodedPacket[3][84] ), .ZN(n6083) );
  NBUFFX2 U6593 ( .INP(n826), .Z(n5851) );
  NBUFFX2 U6594 ( .INP(n5848), .Z(n5850) );
  NBUFFX2 U6595 ( .INP(n5851), .Z(n5849) );
  NBUFFX2 U6596 ( .INP(n5849), .Z(n5848) );
  NBUFFX2 U6597 ( .INP(n5851), .Z(n5853) );
  NBUFFX2 U6598 ( .INP(n826), .Z(n5852) );
  INVX0 U6599 ( .INP(\decodedPacket[3][71] ), .ZN(n6053) );
  INVX0 U6600 ( .INP(\decodedPacket[5][84] ), .ZN(n6237) );
  INVX0 U6601 ( .INP(\decodedPacket[3][72] ), .ZN(n6086) );
  INVX0 U6602 ( .INP(\decodedPacket[5][71] ), .ZN(n6207) );
  NBUFFX2 U6603 ( .INP(n1124), .Z(n5690) );
  INVX0 U6604 ( .INP(\decodedPacket[5][72] ), .ZN(n6240) );
  INVX0 U6605 ( .INP(\decodedPacket[7][84] ), .ZN(n6391) );
  INVX0 U6606 ( .INP(\decodedPacket[7][71] ), .ZN(n6361) );
  INVX0 U6607 ( .INP(\decodedPacket[7][72] ), .ZN(n6394) );
  OAI22X1 U6608 ( .IN1(n5600), .IN2(n1816), .IN3(n6063), .IN4(n5599), .QN(
        n5196) );
  OAI22X1 U6609 ( .IN1(n5600), .IN2(n1792), .IN3(n5854), .IN4(n5614), .QN(
        n5197) );
  INVX0 U6610 ( .INP(\decodedPacket[2][117] ), .ZN(n6063) );
  AND2X1 U6611 ( .IN1(\decodedPacket[2][117] ), .IN2(n5691), .Q(n5198) );
  NAND2X1 U6612 ( .IN1(n5773), .IN2(\decodedPacket[2][117] ), .QN(n4614) );
  NAND2X1 U6613 ( .IN1(n5276), .IN2(\decodedPacket[2][117] ), .QN(n4109) );
  INVX0 U6614 ( .INP(\decodedPacket[2][98] ), .ZN(n5998) );
  INVX0 U6615 ( .INP(\decodedPacket[2][116] ), .ZN(n6062) );
  INVX0 U6616 ( .INP(\decodedPacket[2][91] ), .ZN(n6108) );
  INVX0 U6617 ( .INP(\decodedPacket[2][120] ), .ZN(n6041) );
  INVX0 U6618 ( .INP(\decodedPacket[2][118] ), .ZN(n6066) );
  INVX0 U6619 ( .INP(n1768), .ZN(n5591) );
  INVX0 U6620 ( .INP(n2521), .ZN(\add_177_I3_aco/A[0] ) );
  NBUFFX2 U6621 ( .INP(n1114), .Z(n5766) );
  INVX0 U6622 ( .INP(N2172), .ZN(n5995) );
  NBUFFX4 U6623 ( .INP(n5199), .Z(n5282) );
  NBUFFX4 U6624 ( .INP(n5200), .Z(n5622) );
  INVX0 U6625 ( .INP(N1068), .ZN(n5996) );
  INVX0 U6626 ( .INP(N8580), .ZN(n5992) );
  INVX0 U6627 ( .INP(N4308), .ZN(n5994) );
  INVX0 U6628 ( .INP(n2522), .ZN(\add_177_I3_aco/A[1] ) );
  INVX0 U6629 ( .INP(N6444), .ZN(n5993) );
  NAND2X1 U6630 ( .IN1(\decodedPacket[0][117] ), .IN2(n5586), .QN(n1816) );
  INVX0 U6631 ( .INP(\decodedPacket[4][117] ), .ZN(n6217) );
  NBUFFX2 U6632 ( .INP(decodedVector_o[4]), .Z(n5897) );
  NBUFFX2 U6633 ( .INP(decodedVector_o[4]), .Z(n5898) );
  NBUFFX2 U6634 ( .INP(decodedVector_o[4]), .Z(n5899) );
  NBUFFX2 U6635 ( .INP(decodedVector_o[4]), .Z(n5900) );
  NBUFFX2 U6636 ( .INP(decodedVector_o[4]), .Z(n5901) );
  NBUFFX2 U6637 ( .INP(decodedVector_o[4]), .Z(n5902) );
  NBUFFX2 U6638 ( .INP(decodedVector_o[4]), .Z(n5903) );
  NBUFFX2 U6639 ( .INP(decodedVector_o[4]), .Z(n5904) );
  NBUFFX2 U6640 ( .INP(decodedVector_o[4]), .Z(n5905) );
  NBUFFX2 U6641 ( .INP(decodedVector_o[4]), .Z(n5906) );
  NBUFFX2 U6642 ( .INP(decodedVector_o[5]), .Z(n5907) );
  NBUFFX2 U6643 ( .INP(decodedVector_o[5]), .Z(n5908) );
  NBUFFX2 U6644 ( .INP(decodedVector_o[5]), .Z(n5909) );
  NBUFFX2 U6645 ( .INP(decodedVector_o[5]), .Z(n5910) );
  NBUFFX2 U6646 ( .INP(decodedVector_o[5]), .Z(n5911) );
  NBUFFX2 U6647 ( .INP(decodedVector_o[5]), .Z(n5912) );
  NBUFFX2 U6648 ( .INP(decodedVector_o[5]), .Z(n5913) );
  NBUFFX2 U6649 ( .INP(decodedVector_o[5]), .Z(n5914) );
  NBUFFX2 U6650 ( .INP(decodedVector_o[5]), .Z(n5915) );
  NBUFFX2 U6651 ( .INP(decodedVector_o[5]), .Z(n5916) );
  NBUFFX2 U6652 ( .INP(decodedVector_o[6]), .Z(n5917) );
  NBUFFX2 U6653 ( .INP(decodedVector_o[6]), .Z(n5918) );
  NBUFFX2 U6654 ( .INP(decodedVector_o[6]), .Z(n5919) );
  NBUFFX2 U6655 ( .INP(decodedVector_o[6]), .Z(n5920) );
  NBUFFX2 U6656 ( .INP(decodedVector_o[6]), .Z(n5921) );
  NBUFFX2 U6657 ( .INP(decodedVector_o[6]), .Z(n5922) );
  NBUFFX2 U6658 ( .INP(decodedVector_o[6]), .Z(n5923) );
  NBUFFX2 U6659 ( .INP(decodedVector_o[6]), .Z(n5924) );
  NBUFFX2 U6660 ( .INP(decodedVector_o[6]), .Z(n5925) );
  NBUFFX2 U6661 ( .INP(decodedVector_o[6]), .Z(n5926) );
  NBUFFX2 U6662 ( .INP(decodedVector_o[7]), .Z(n5927) );
  NBUFFX2 U6663 ( .INP(decodedVector_o[7]), .Z(n5928) );
  NBUFFX2 U6664 ( .INP(decodedVector_o[7]), .Z(n5929) );
  NBUFFX2 U6665 ( .INP(decodedVector_o[7]), .Z(n5930) );
  NBUFFX2 U6666 ( .INP(decodedVector_o[7]), .Z(n5931) );
  NBUFFX2 U6667 ( .INP(decodedVector_o[7]), .Z(n5932) );
  NBUFFX2 U6668 ( .INP(decodedVector_o[7]), .Z(n5933) );
  NBUFFX2 U6669 ( .INP(decodedVector_o[7]), .Z(n5934) );
  NBUFFX2 U6670 ( .INP(decodedVector_o[7]), .Z(n5935) );
  NBUFFX2 U6671 ( .INP(decodedVector_o[7]), .Z(n5936) );
  NBUFFX2 U6672 ( .INP(decodedVector_o[0]), .Z(n5857) );
  NBUFFX2 U6673 ( .INP(decodedVector_o[0]), .Z(n5858) );
  NBUFFX2 U6674 ( .INP(decodedVector_o[0]), .Z(n5859) );
  NBUFFX2 U6675 ( .INP(decodedVector_o[0]), .Z(n5860) );
  NBUFFX2 U6676 ( .INP(decodedVector_o[0]), .Z(n5861) );
  NBUFFX2 U6677 ( .INP(decodedVector_o[0]), .Z(n5862) );
  NBUFFX2 U6678 ( .INP(decodedVector_o[0]), .Z(n5863) );
  NBUFFX2 U6679 ( .INP(decodedVector_o[0]), .Z(n5864) );
  NBUFFX2 U6680 ( .INP(decodedVector_o[0]), .Z(n5865) );
  NBUFFX2 U6681 ( .INP(decodedVector_o[0]), .Z(n5866) );
  NBUFFX2 U6682 ( .INP(decodedVector_o[2]), .Z(n5877) );
  NBUFFX2 U6683 ( .INP(decodedVector_o[2]), .Z(n5878) );
  NBUFFX2 U6684 ( .INP(decodedVector_o[2]), .Z(n5879) );
  NBUFFX2 U6685 ( .INP(decodedVector_o[2]), .Z(n5880) );
  NBUFFX2 U6686 ( .INP(decodedVector_o[2]), .Z(n5881) );
  NBUFFX2 U6687 ( .INP(decodedVector_o[2]), .Z(n5882) );
  NBUFFX2 U6688 ( .INP(decodedVector_o[2]), .Z(n5883) );
  NBUFFX2 U6689 ( .INP(decodedVector_o[2]), .Z(n5884) );
  NBUFFX2 U6690 ( .INP(decodedVector_o[2]), .Z(n5885) );
  NBUFFX2 U6691 ( .INP(decodedVector_o[2]), .Z(n5886) );
  NBUFFX2 U6692 ( .INP(n1763), .Z(n5628) );
  NBUFFX2 U6693 ( .INP(n1763), .Z(n5629) );
  NBUFFX2 U6694 ( .INP(n1763), .Z(n5630) );
  NBUFFX2 U6695 ( .INP(n1763), .Z(n5631) );
  NBUFFX2 U6696 ( .INP(n1763), .Z(n5632) );
  NBUFFX2 U6697 ( .INP(n1763), .Z(n5633) );
  NBUFFX2 U6698 ( .INP(n1763), .Z(n5634) );
  NBUFFX2 U6699 ( .INP(n1763), .Z(n5635) );
  INVX0 U6700 ( .INP(\decodedPacket[6][117] ), .ZN(n6371) );
  NBUFFX2 U6701 ( .INP(n1114), .Z(n5771) );
  INVX0 U6702 ( .INP(\decodedPacket[4][116] ), .ZN(n6216) );
  INVX0 U6703 ( .INP(\decodedPacket[6][116] ), .ZN(n6370) );
  INVX0 U6704 ( .INP(\decodedPacket[4][91] ), .ZN(n6262) );
  INVX0 U6705 ( .INP(\decodedPacket[6][91] ), .ZN(n6416) );
  NBUFFX2 U6706 ( .INP(n1114), .Z(n5770) );
  INVX0 U6707 ( .INP(\decodedPacket[4][120] ), .ZN(n6195) );
  INVX0 U6708 ( .INP(\decodedPacket[6][120] ), .ZN(n6349) );
  NBUFFX2 U6709 ( .INP(n1114), .Z(n5769) );
  NBUFFX2 U6710 ( .INP(n1114), .Z(n5768) );
  NBUFFX2 U6711 ( .INP(n1114), .Z(n5767) );
  NBUFFX2 U6712 ( .INP(n1763), .Z(n5636) );
  NBUFFX2 U6713 ( .INP(n1767), .Z(n5597) );
  NBUFFX2 U6714 ( .INP(n1767), .Z(n5598) );
  NBUFFX2 U6715 ( .INP(n1767), .Z(n5599) );
  NBUFFX2 U6716 ( .INP(n1114), .Z(n5772) );
  NBUFFX2 U6717 ( .INP(n3680), .Z(n5397) );
  NBUFFX2 U6718 ( .INP(n3296), .Z(n5456) );
  NBUFFX2 U6719 ( .INP(n2912), .Z(n5515) );
  NBUFFX2 U6720 ( .INP(n2523), .Z(n5573) );
  NBUFFX2 U6721 ( .INP(n2523), .Z(n5574) );
  NBUFFX2 U6722 ( .INP(n832), .Z(n5789) );
  NBUFFX2 U6723 ( .INP(n832), .Z(n5788) );
  NBUFFX2 U6724 ( .INP(n832), .Z(n5787) );
  NBUFFX2 U6725 ( .INP(n828), .Z(n5825) );
  NBUFFX2 U6726 ( .INP(n828), .Z(n5824) );
  NBUFFX2 U6727 ( .INP(n828), .Z(n5823) );
  NBUFFX2 U6728 ( .INP(n828), .Z(n5822) );
  NBUFFX2 U6729 ( .INP(n3680), .Z(n5398) );
  NBUFFX2 U6730 ( .INP(n3296), .Z(n5457) );
  NBUFFX2 U6731 ( .INP(n2912), .Z(n5516) );
  NBUFFX2 U6732 ( .INP(n2523), .Z(n5575) );
  INVX0 U6733 ( .INP(n1768), .ZN(n5595) );
  INVX0 U6734 ( .INP(n1768), .ZN(n5594) );
  INVX0 U6735 ( .INP(n1768), .ZN(n5593) );
  INVX0 U6736 ( .INP(n1768), .ZN(n5592) );
  NBUFFX4 U6737 ( .INP(n5200), .Z(n5623) );
  NBUFFX2 U6738 ( .INP(n5199), .Z(n5283) );
  INVX0 U6739 ( .INP(\decodedPacket[2][107] ), .ZN(n6054) );
  INVX0 U6740 ( .INP(\decodedPacket[2][108] ), .ZN(n6055) );
  INVX0 U6741 ( .INP(\decodedPacket[2][109] ), .ZN(n6056) );
  INVX0 U6742 ( .INP(\decodedPacket[2][110] ), .ZN(n6057) );
  INVX0 U6743 ( .INP(\decodedPacket[2][111] ), .ZN(n6058) );
  INVX0 U6744 ( .INP(\decodedPacket[2][85] ), .ZN(n6046) );
  INVX0 U6745 ( .INP(\decodedPacket[2][86] ), .ZN(n6047) );
  INVX0 U6746 ( .INP(\decodedPacket[2][87] ), .ZN(n6048) );
  INVX0 U6747 ( .INP(\decodedPacket[2][88] ), .ZN(n6049) );
  INVX0 U6748 ( .INP(\decodedPacket[2][89] ), .ZN(n6050) );
  INVX0 U6749 ( .INP(\decodedPacket[2][90] ), .ZN(n6051) );
  INVX0 U6750 ( .INP(n1768), .ZN(n5596) );
  INVX0 U6751 ( .INP(\decodedPacket[2][73] ), .ZN(n6097) );
  INVX0 U6752 ( .INP(\decodedPacket[2][74] ), .ZN(n6096) );
  INVX0 U6753 ( .INP(\decodedPacket[2][75] ), .ZN(n6095) );
  INVX0 U6754 ( .INP(\decodedPacket[2][76] ), .ZN(n6094) );
  INVX0 U6755 ( .INP(\decodedPacket[2][83] ), .ZN(n6107) );
  INVX0 U6756 ( .INP(\decodedPacket[2][94] ), .ZN(n6111) );
  INVX0 U6757 ( .INP(\decodedPacket[2][95] ), .ZN(n6112) );
  INVX0 U6758 ( .INP(\decodedPacket[2][92] ), .ZN(n6109) );
  INVX0 U6759 ( .INP(\decodedPacket[2][96] ), .ZN(n6113) );
  INVX0 U6760 ( .INP(\decodedPacket[2][78] ), .ZN(n6102) );
  INVX0 U6761 ( .INP(\decodedPacket[2][93] ), .ZN(n6110) );
  INVX0 U6762 ( .INP(\decodedPacket[2][71] ), .ZN(n6052) );
  NAND2X1 U6763 ( .IN1(decodedPacketValid[1]), .IN2(n5997), .QN(n1768) );
  NOR2X0 U6764 ( .IN1(n5401), .IN2(n5351), .QN(n4063) );
  NOR2X0 U6765 ( .IN1(n5460), .IN2(n5410), .QN(n3679) );
  NOR2X0 U6766 ( .IN1(n5519), .IN2(n5469), .QN(n3295) );
  NOR2X0 U6767 ( .IN1(n5578), .IN2(n5528), .QN(n2906) );
  INVX0 U6768 ( .INP(N389), .ZN(n5997) );
  NOR4X0 U6769 ( .IN1(decodedPacketValid[1]), .IN2(N389), .IN3(n5673), .IN4(
        n5600), .QN(n2520) );
  NOR2X0 U6770 ( .IN1(n5622), .IN2(n5624), .QN(n2519) );
  AND4X1 U6771 ( .IN1(n5986), .IN2(decodedPacketValid[3]), .IN3(N1069), .IN4(
        N1068), .Q(n5199) );
  AND4X1 U6772 ( .IN1(n5986), .IN2(decodedPacketValid[3]), .IN3(n5996), .IN4(
        n5991), .Q(n5200) );
  NAND2X1 U6773 ( .IN1(decodedPacketValid[2]), .IN2(\add_177_I3_aco/A[1] ), 
        .QN(n4691) );
  AND4X1 U6774 ( .IN1(n5986), .IN2(decodedPacketValid[3]), .IN3(N1068), .IN4(
        n5991), .Q(n5201) );
  NAND2X1 U6775 ( .IN1(decodedPacketValid[1]), .IN2(N389), .QN(n2522) );
  NAND2X1 U6776 ( .IN1(decodedPacketValid[2]), .IN2(\add_177_I3_aco/A[0] ), 
        .QN(n1124) );
  NAND3X0 U6777 ( .IN1(n2521), .IN2(n2522), .IN3(decodedPacketValid[2]), .QN(
        n1767) );
  NOR2X0 U6778 ( .IN1(n2483), .IN2(n5673), .QN(N9674) );
  NAND2X1 U6779 ( .IN1(n5639), .IN2(n5044), .QN(n2484) );
  NOR2X0 U6780 ( .IN1(n2477), .IN2(n5673), .QN(N9675) );
  NAND2X1 U6781 ( .IN1(n5639), .IN2(n5045), .QN(n2478) );
  NOR2X0 U6782 ( .IN1(n2471), .IN2(n5673), .QN(N9676) );
  NAND2X1 U6783 ( .IN1(n5639), .IN2(n5046), .QN(n2472) );
  NOR2X0 U6784 ( .IN1(n2465), .IN2(n5673), .QN(N9677) );
  NAND2X1 U6785 ( .IN1(n5639), .IN2(n5047), .QN(n2466) );
  NOR2X0 U6786 ( .IN1(n2459), .IN2(n5673), .QN(N9678) );
  NAND2X1 U6787 ( .IN1(n5639), .IN2(n5048), .QN(n2460) );
  NOR2X0 U6788 ( .IN1(n2453), .IN2(n5673), .QN(N9679) );
  NAND2X1 U6789 ( .IN1(n5639), .IN2(n5049), .QN(n2454) );
  NOR2X0 U6790 ( .IN1(n2447), .IN2(n5673), .QN(N9680) );
  NAND2X1 U6791 ( .IN1(n5639), .IN2(n5050), .QN(n2448) );
  NOR2X0 U6792 ( .IN1(n2441), .IN2(n5673), .QN(N9681) );
  NAND2X1 U6793 ( .IN1(n5639), .IN2(n5051), .QN(n2442) );
  NOR2X0 U6794 ( .IN1(n2435), .IN2(n5673), .QN(N9682) );
  NAND2X1 U6795 ( .IN1(n5639), .IN2(n5052), .QN(n2436) );
  NOR2X0 U6796 ( .IN1(n2429), .IN2(n5673), .QN(N9683) );
  NAND2X1 U6797 ( .IN1(n5639), .IN2(n5053), .QN(n2430) );
  NOR2X0 U6798 ( .IN1(n1720), .IN2(n5763), .QN(N9803) );
  NAND2X1 U6799 ( .IN1(n5729), .IN2(n5157), .QN(n1721) );
  NOR2X0 U6800 ( .IN1(n1715), .IN2(n5763), .QN(N9804) );
  NAND2X1 U6801 ( .IN1(n5729), .IN2(n5158), .QN(n1716) );
  NOR2X0 U6802 ( .IN1(n1710), .IN2(n5763), .QN(N9805) );
  NAND2X1 U6803 ( .IN1(n5729), .IN2(n5159), .QN(n1711) );
  NOR2X0 U6804 ( .IN1(n1705), .IN2(n5763), .QN(N9806) );
  NAND2X1 U6805 ( .IN1(n5729), .IN2(n5160), .QN(n1706) );
  NOR2X0 U6806 ( .IN1(n1700), .IN2(n5763), .QN(N9807) );
  NAND2X1 U6807 ( .IN1(n5729), .IN2(n5161), .QN(n1701) );
  NOR2X0 U6808 ( .IN1(n1695), .IN2(n5763), .QN(N9808) );
  NAND2X1 U6809 ( .IN1(n5729), .IN2(n5162), .QN(n1696) );
  NOR2X0 U6810 ( .IN1(n1690), .IN2(n5763), .QN(N9809) );
  NAND2X1 U6811 ( .IN1(n5729), .IN2(n5163), .QN(n1691) );
  NOR2X0 U6812 ( .IN1(n1685), .IN2(n5763), .QN(N9810) );
  NAND2X1 U6813 ( .IN1(n5729), .IN2(n5062), .QN(n1686) );
  NOR2X0 U6814 ( .IN1(n1680), .IN2(n5763), .QN(N9811) );
  NAND2X1 U6815 ( .IN1(n5729), .IN2(n5063), .QN(n1681) );
  NOR2X0 U6816 ( .IN1(n1675), .IN2(n5763), .QN(N9812) );
  NAND2X1 U6817 ( .IN1(n5729), .IN2(n5064), .QN(n1676) );
  NOR2X0 U6818 ( .IN1(n4554), .IN2(n5340), .QN(N10063) );
  NAND2X1 U6819 ( .IN1(n5306), .IN2(n5091), .QN(n4555) );
  NOR2X0 U6820 ( .IN1(n4550), .IN2(n5340), .QN(N10064) );
  NAND2X1 U6821 ( .IN1(n5306), .IN2(n5092), .QN(n4551) );
  NOR2X0 U6822 ( .IN1(n4546), .IN2(n5340), .QN(N10065) );
  NAND2X1 U6823 ( .IN1(n5306), .IN2(n5093), .QN(n4547) );
  NOR2X0 U6824 ( .IN1(n4542), .IN2(n5340), .QN(N10066) );
  NAND2X1 U6825 ( .IN1(n5306), .IN2(n5094), .QN(n4543) );
  NOR2X0 U6826 ( .IN1(n4538), .IN2(n5340), .QN(N10067) );
  NAND2X1 U6827 ( .IN1(n5306), .IN2(n5095), .QN(n4539) );
  NOR2X0 U6828 ( .IN1(n4534), .IN2(n5340), .QN(N10068) );
  NAND2X1 U6829 ( .IN1(n5306), .IN2(n5096), .QN(n4535) );
  NOR2X0 U6830 ( .IN1(n4530), .IN2(n5340), .QN(N10069) );
  NAND2X1 U6831 ( .IN1(n5306), .IN2(n5097), .QN(n4531) );
  NOR2X0 U6832 ( .IN1(n4526), .IN2(n5340), .QN(N10070) );
  NAND2X1 U6833 ( .IN1(n5306), .IN2(n5098), .QN(n4527) );
  NOR2X0 U6834 ( .IN1(n4522), .IN2(n5340), .QN(N10071) );
  NAND2X1 U6835 ( .IN1(n5306), .IN2(n5099), .QN(n4523) );
  NOR2X0 U6836 ( .IN1(n4518), .IN2(n5340), .QN(N10072) );
  NAND2X1 U6837 ( .IN1(n5306), .IN2(n5100), .QN(n4519) );
  NOR2X0 U6838 ( .IN1(n4044), .IN2(n5401), .QN(N10193) );
  NAND2X1 U6839 ( .IN1(n5365), .IN2(n5164), .QN(n4045) );
  NOR2X0 U6840 ( .IN1(n4041), .IN2(n5401), .QN(N10194) );
  NAND2X1 U6841 ( .IN1(n5365), .IN2(n5165), .QN(n4042) );
  NOR2X0 U6842 ( .IN1(n4038), .IN2(n5401), .QN(N10195) );
  NAND2X1 U6843 ( .IN1(n5365), .IN2(n5166), .QN(n4039) );
  NOR2X0 U6844 ( .IN1(n4035), .IN2(n5401), .QN(N10196) );
  NAND2X1 U6845 ( .IN1(n5365), .IN2(n5167), .QN(n4036) );
  NOR2X0 U6846 ( .IN1(n4032), .IN2(n5401), .QN(N10197) );
  NAND2X1 U6847 ( .IN1(n5365), .IN2(n5168), .QN(n4033) );
  NOR2X0 U6848 ( .IN1(n4029), .IN2(n5401), .QN(N10198) );
  NAND2X1 U6849 ( .IN1(n5365), .IN2(n5169), .QN(n4030) );
  NOR2X0 U6850 ( .IN1(n4026), .IN2(n5401), .QN(N10199) );
  NAND2X1 U6851 ( .IN1(n5365), .IN2(n4945), .QN(n4027) );
  NOR2X0 U6852 ( .IN1(n4023), .IN2(n5401), .QN(N10200) );
  NAND2X1 U6853 ( .IN1(n5365), .IN2(n5170), .QN(n4024) );
  NOR2X0 U6854 ( .IN1(n4020), .IN2(n5401), .QN(N10201) );
  NAND2X1 U6855 ( .IN1(n5365), .IN2(n4946), .QN(n4021) );
  NOR2X0 U6856 ( .IN1(n4017), .IN2(n5401), .QN(N10202) );
  NAND2X1 U6857 ( .IN1(n5365), .IN2(n4947), .QN(n4018) );
  NOR2X0 U6858 ( .IN1(n3660), .IN2(n5460), .QN(N10323) );
  NAND2X1 U6859 ( .IN1(n5424), .IN2(n5171), .QN(n3661) );
  NOR2X0 U6860 ( .IN1(n3657), .IN2(n5460), .QN(N10324) );
  NAND2X1 U6861 ( .IN1(n5424), .IN2(n5172), .QN(n3658) );
  NOR2X0 U6862 ( .IN1(n3654), .IN2(n5460), .QN(N10325) );
  NAND2X1 U6863 ( .IN1(n5424), .IN2(n5173), .QN(n3655) );
  NOR2X0 U6864 ( .IN1(n3651), .IN2(n5460), .QN(N10326) );
  NAND2X1 U6865 ( .IN1(n5424), .IN2(n5174), .QN(n3652) );
  NOR2X0 U6866 ( .IN1(n3648), .IN2(n5460), .QN(N10327) );
  NAND2X1 U6867 ( .IN1(n5424), .IN2(n5175), .QN(n3649) );
  NOR2X0 U6868 ( .IN1(n3645), .IN2(n5460), .QN(N10328) );
  NAND2X1 U6869 ( .IN1(n5424), .IN2(n5176), .QN(n3646) );
  NOR2X0 U6870 ( .IN1(n3642), .IN2(n5460), .QN(N10329) );
  NAND2X1 U6871 ( .IN1(n5424), .IN2(n4948), .QN(n3643) );
  NOR2X0 U6872 ( .IN1(n3639), .IN2(n5460), .QN(N10330) );
  NAND2X1 U6873 ( .IN1(n5424), .IN2(n5177), .QN(n3640) );
  NOR2X0 U6874 ( .IN1(n3636), .IN2(n5460), .QN(N10331) );
  NAND2X1 U6875 ( .IN1(n5424), .IN2(n4949), .QN(n3637) );
  NOR2X0 U6876 ( .IN1(n3633), .IN2(n5460), .QN(N10332) );
  NAND2X1 U6877 ( .IN1(n5424), .IN2(n4950), .QN(n3634) );
  NOR2X0 U6878 ( .IN1(n3276), .IN2(n5519), .QN(N10453) );
  NAND2X1 U6879 ( .IN1(n5483), .IN2(n5178), .QN(n3277) );
  NOR2X0 U6880 ( .IN1(n3273), .IN2(n5519), .QN(N10454) );
  NAND2X1 U6881 ( .IN1(n5483), .IN2(n5179), .QN(n3274) );
  NOR2X0 U6882 ( .IN1(n3270), .IN2(n5519), .QN(N10455) );
  NAND2X1 U6883 ( .IN1(n5483), .IN2(n5180), .QN(n3271) );
  NOR2X0 U6884 ( .IN1(n3267), .IN2(n5519), .QN(N10456) );
  NAND2X1 U6885 ( .IN1(n5483), .IN2(n5181), .QN(n3268) );
  NOR2X0 U6886 ( .IN1(n3264), .IN2(n5519), .QN(N10457) );
  NAND2X1 U6887 ( .IN1(n5483), .IN2(n5182), .QN(n3265) );
  NOR2X0 U6888 ( .IN1(n3261), .IN2(n5519), .QN(N10458) );
  NAND2X1 U6889 ( .IN1(n5483), .IN2(n5183), .QN(n3262) );
  NOR2X0 U6890 ( .IN1(n3258), .IN2(n5519), .QN(N10459) );
  NAND2X1 U6891 ( .IN1(n5483), .IN2(n4951), .QN(n3259) );
  NOR2X0 U6892 ( .IN1(n3255), .IN2(n5519), .QN(N10460) );
  NAND2X1 U6893 ( .IN1(n5483), .IN2(n5184), .QN(n3256) );
  NOR2X0 U6894 ( .IN1(n3252), .IN2(n5519), .QN(N10461) );
  NAND2X1 U6895 ( .IN1(n5483), .IN2(n4952), .QN(n3253) );
  NOR2X0 U6896 ( .IN1(n3249), .IN2(n5519), .QN(N10462) );
  NAND2X1 U6897 ( .IN1(n5483), .IN2(n4953), .QN(n3250) );
  NOR2X0 U6898 ( .IN1(n2887), .IN2(n5578), .QN(N10583) );
  NAND2X1 U6899 ( .IN1(n5541), .IN2(n5185), .QN(n2888) );
  NOR2X0 U6900 ( .IN1(n2884), .IN2(n5578), .QN(N10584) );
  NAND2X1 U6901 ( .IN1(n5541), .IN2(n5186), .QN(n2885) );
  NOR2X0 U6902 ( .IN1(n2881), .IN2(n5578), .QN(N10585) );
  NAND2X1 U6903 ( .IN1(n5541), .IN2(n5187), .QN(n2882) );
  NOR2X0 U6904 ( .IN1(n2878), .IN2(n5578), .QN(N10586) );
  NAND2X1 U6905 ( .IN1(n5541), .IN2(n5188), .QN(n2879) );
  NOR2X0 U6906 ( .IN1(n2875), .IN2(n5578), .QN(N10587) );
  NAND2X1 U6907 ( .IN1(n5541), .IN2(n5189), .QN(n2876) );
  NOR2X0 U6908 ( .IN1(n2872), .IN2(n5578), .QN(N10588) );
  NAND2X1 U6909 ( .IN1(n5541), .IN2(n5190), .QN(n2873) );
  NOR2X0 U6910 ( .IN1(n2869), .IN2(n5578), .QN(N10589) );
  NAND2X1 U6911 ( .IN1(n5541), .IN2(n4920), .QN(n2870) );
  NOR2X0 U6912 ( .IN1(n2866), .IN2(n5578), .QN(N10590) );
  NAND2X1 U6913 ( .IN1(n5541), .IN2(n5191), .QN(n2867) );
  NOR2X0 U6914 ( .IN1(n2863), .IN2(n5578), .QN(N10591) );
  NAND2X1 U6915 ( .IN1(n5541), .IN2(n4921), .QN(n2864) );
  NOR2X0 U6916 ( .IN1(n2860), .IN2(n5578), .QN(N10592) );
  NAND2X1 U6917 ( .IN1(n5541), .IN2(n4922), .QN(n2861) );
  NOR2X0 U6918 ( .IN1(n1090), .IN2(n5845), .QN(N9933) );
  NAND2X1 U6919 ( .IN1(n5810), .IN2(n5125), .QN(n1091) );
  NOR2X0 U6920 ( .IN1(n1086), .IN2(n5845), .QN(N9934) );
  NAND2X1 U6921 ( .IN1(n5810), .IN2(n5126), .QN(n1087) );
  NOR2X0 U6922 ( .IN1(n1082), .IN2(n5845), .QN(N9935) );
  NAND2X1 U6923 ( .IN1(n5810), .IN2(n5127), .QN(n1083) );
  NOR2X0 U6924 ( .IN1(n1078), .IN2(n5845), .QN(N9936) );
  NAND2X1 U6925 ( .IN1(n5810), .IN2(n5128), .QN(n1079) );
  NOR2X0 U6926 ( .IN1(n1074), .IN2(n5845), .QN(N9937) );
  NAND2X1 U6927 ( .IN1(n5810), .IN2(n5129), .QN(n1075) );
  NOR2X0 U6928 ( .IN1(n1070), .IN2(n5845), .QN(N9938) );
  NAND2X1 U6929 ( .IN1(n5810), .IN2(n5130), .QN(n1071) );
  NOR2X0 U6930 ( .IN1(n1066), .IN2(n5845), .QN(N9939) );
  NAND2X1 U6931 ( .IN1(n5810), .IN2(n5131), .QN(n1067) );
  NOR2X0 U6932 ( .IN1(n1062), .IN2(n5845), .QN(N9940) );
  NAND2X1 U6933 ( .IN1(n5810), .IN2(n5132), .QN(n1063) );
  NOR2X0 U6934 ( .IN1(n1058), .IN2(n5845), .QN(N9941) );
  NAND2X1 U6935 ( .IN1(n5810), .IN2(n5133), .QN(n1059) );
  NOR2X0 U6936 ( .IN1(n1054), .IN2(n5845), .QN(N9942) );
  NAND2X1 U6937 ( .IN1(n5810), .IN2(n5134), .QN(n1055) );
  NOR2X0 U6938 ( .IN1(n1670), .IN2(n5762), .QN(N9813) );
  NAND2X1 U6939 ( .IN1(n5728), .IN2(n5065), .QN(n1671) );
  NOR2X0 U6940 ( .IN1(n1665), .IN2(n5762), .QN(N9814) );
  NAND2X1 U6941 ( .IN1(n5728), .IN2(n5066), .QN(n1666) );
  NOR2X0 U6942 ( .IN1(n1660), .IN2(n5762), .QN(N9815) );
  NAND2X1 U6943 ( .IN1(n5728), .IN2(n5067), .QN(n1661) );
  NOR2X0 U6944 ( .IN1(n1655), .IN2(n5762), .QN(N9816) );
  NAND2X1 U6945 ( .IN1(n5728), .IN2(n5068), .QN(n1656) );
  NOR2X0 U6946 ( .IN1(n1650), .IN2(n5762), .QN(N9817) );
  NAND2X1 U6947 ( .IN1(n5728), .IN2(n5069), .QN(n1651) );
  NOR2X0 U6948 ( .IN1(n1645), .IN2(n5762), .QN(N9818) );
  NAND2X1 U6949 ( .IN1(n5728), .IN2(n5070), .QN(n1646) );
  NOR2X0 U6950 ( .IN1(n1640), .IN2(n5762), .QN(N9819) );
  NAND2X1 U6951 ( .IN1(n5728), .IN2(n5071), .QN(n1641) );
  NOR2X0 U6952 ( .IN1(n1635), .IN2(n5762), .QN(N9820) );
  NAND2X1 U6953 ( .IN1(n5728), .IN2(n5072), .QN(n1636) );
  NOR2X0 U6954 ( .IN1(n1630), .IN2(n5762), .QN(N9821) );
  NAND2X1 U6955 ( .IN1(n5728), .IN2(n5073), .QN(n1631) );
  NOR2X0 U6956 ( .IN1(n1625), .IN2(n5762), .QN(N9822) );
  NAND2X1 U6957 ( .IN1(n5728), .IN2(n5074), .QN(n1626) );
  NOR2X0 U6958 ( .IN1(n1620), .IN2(n5762), .QN(N9823) );
  NAND2X1 U6959 ( .IN1(n5728), .IN2(n5075), .QN(n1621) );
  NOR2X0 U6960 ( .IN1(n1615), .IN2(n5762), .QN(N9824) );
  NAND2X1 U6961 ( .IN1(n5728), .IN2(n5076), .QN(n1616) );
  NOR2X0 U6962 ( .IN1(n1610), .IN2(n5761), .QN(N9825) );
  NAND2X1 U6963 ( .IN1(n5727), .IN2(n5077), .QN(n1611) );
  NOR2X0 U6964 ( .IN1(n1605), .IN2(n5761), .QN(N9826) );
  NAND2X1 U6965 ( .IN1(n5727), .IN2(n5078), .QN(n1606) );
  NOR2X0 U6966 ( .IN1(n1600), .IN2(n5761), .QN(N9827) );
  NAND2X1 U6967 ( .IN1(n5727), .IN2(n5079), .QN(n1601) );
  NOR2X0 U6968 ( .IN1(n1595), .IN2(n5761), .QN(N9828) );
  NAND2X1 U6969 ( .IN1(n5727), .IN2(n5080), .QN(n1596) );
  NOR2X0 U6970 ( .IN1(n1590), .IN2(n5761), .QN(N9829) );
  NAND2X1 U6971 ( .IN1(n5727), .IN2(n5081), .QN(n1591) );
  NOR2X0 U6972 ( .IN1(n1585), .IN2(n5761), .QN(N9830) );
  NAND2X1 U6973 ( .IN1(n5727), .IN2(n5082), .QN(n1586) );
  NOR2X0 U6974 ( .IN1(n1580), .IN2(n5761), .QN(N9831) );
  NAND2X1 U6975 ( .IN1(n5727), .IN2(n5083), .QN(n1581) );
  NOR2X0 U6976 ( .IN1(n1575), .IN2(n5761), .QN(N9832) );
  NAND2X1 U6977 ( .IN1(n5727), .IN2(n5084), .QN(n1576) );
  NOR2X0 U6978 ( .IN1(n1570), .IN2(n5761), .QN(N9833) );
  NAND2X1 U6979 ( .IN1(n5727), .IN2(n5085), .QN(n1571) );
  NOR2X0 U6980 ( .IN1(n1565), .IN2(n5761), .QN(N9834) );
  NAND2X1 U6981 ( .IN1(n5727), .IN2(n5086), .QN(n1566) );
  NOR2X0 U6982 ( .IN1(n3978), .IN2(n5399), .QN(N10215) );
  NAND2X1 U6983 ( .IN1(n5363), .IN2(n4995), .QN(n3979) );
  NOR2X0 U6984 ( .IN1(n3975), .IN2(n5399), .QN(N10216) );
  NAND2X1 U6985 ( .IN1(n5363), .IN2(n4996), .QN(n3976) );
  NOR2X0 U6986 ( .IN1(n3972), .IN2(n5399), .QN(N10217) );
  NAND2X1 U6987 ( .IN1(n5363), .IN2(n4997), .QN(n3973) );
  NOR2X0 U6988 ( .IN1(n3969), .IN2(n5399), .QN(N10218) );
  NAND2X1 U6989 ( .IN1(n5363), .IN2(n4998), .QN(n3970) );
  NOR2X0 U6990 ( .IN1(n3966), .IN2(n5399), .QN(N10219) );
  NAND2X1 U6991 ( .IN1(n5363), .IN2(n4999), .QN(n3967) );
  NOR2X0 U6992 ( .IN1(n3963), .IN2(n5399), .QN(N10220) );
  NAND2X1 U6993 ( .IN1(n5363), .IN2(n5000), .QN(n3964) );
  NOR2X0 U6994 ( .IN1(n3960), .IN2(n5399), .QN(N10221) );
  NAND2X1 U6995 ( .IN1(n5363), .IN2(n5001), .QN(n3961) );
  NOR2X0 U6996 ( .IN1(n3957), .IN2(n5399), .QN(N10222) );
  NAND2X1 U6997 ( .IN1(n5363), .IN2(n5002), .QN(n3958) );
  NOR2X0 U6998 ( .IN1(n3954), .IN2(n5399), .QN(N10223) );
  NAND2X1 U6999 ( .IN1(n5363), .IN2(n5003), .QN(n3955) );
  NOR2X0 U7000 ( .IN1(n3951), .IN2(n5399), .QN(N10224) );
  NAND2X1 U7001 ( .IN1(n5363), .IN2(n5004), .QN(n3952) );
  NOR2X0 U7002 ( .IN1(n3594), .IN2(n5458), .QN(N10345) );
  NAND2X1 U7003 ( .IN1(n5422), .IN2(n5005), .QN(n3595) );
  NOR2X0 U7004 ( .IN1(n3591), .IN2(n5458), .QN(N10346) );
  NAND2X1 U7005 ( .IN1(n5422), .IN2(n5006), .QN(n3592) );
  NOR2X0 U7006 ( .IN1(n3588), .IN2(n5458), .QN(N10347) );
  NAND2X1 U7007 ( .IN1(n5422), .IN2(n5007), .QN(n3589) );
  NOR2X0 U7008 ( .IN1(n3585), .IN2(n5458), .QN(N10348) );
  NAND2X1 U7009 ( .IN1(n5422), .IN2(n5008), .QN(n3586) );
  NOR2X0 U7010 ( .IN1(n3582), .IN2(n5458), .QN(N10349) );
  NAND2X1 U7011 ( .IN1(n5422), .IN2(n5009), .QN(n3583) );
  NOR2X0 U7012 ( .IN1(n3579), .IN2(n5458), .QN(N10350) );
  NAND2X1 U7013 ( .IN1(n5422), .IN2(n5010), .QN(n3580) );
  NOR2X0 U7014 ( .IN1(n3576), .IN2(n5458), .QN(N10351) );
  NAND2X1 U7015 ( .IN1(n5422), .IN2(n5011), .QN(n3577) );
  NOR2X0 U7016 ( .IN1(n3573), .IN2(n5458), .QN(N10352) );
  NAND2X1 U7017 ( .IN1(n5422), .IN2(n5012), .QN(n3574) );
  NOR2X0 U7018 ( .IN1(n3570), .IN2(n5458), .QN(N10353) );
  NAND2X1 U7019 ( .IN1(n5422), .IN2(n5013), .QN(n3571) );
  NOR2X0 U7020 ( .IN1(n3567), .IN2(n5458), .QN(N10354) );
  NAND2X1 U7021 ( .IN1(n5422), .IN2(n5014), .QN(n3568) );
  NOR2X0 U7022 ( .IN1(n3210), .IN2(n5517), .QN(N10475) );
  NAND2X1 U7023 ( .IN1(n5481), .IN2(n5015), .QN(n3211) );
  NOR2X0 U7024 ( .IN1(n3207), .IN2(n5517), .QN(N10476) );
  NAND2X1 U7025 ( .IN1(n5481), .IN2(n5016), .QN(n3208) );
  NOR2X0 U7026 ( .IN1(n3204), .IN2(n5517), .QN(N10477) );
  NAND2X1 U7027 ( .IN1(n5481), .IN2(n5017), .QN(n3205) );
  NOR2X0 U7028 ( .IN1(n3201), .IN2(n5517), .QN(N10478) );
  NAND2X1 U7029 ( .IN1(n5481), .IN2(n5018), .QN(n3202) );
  NOR2X0 U7030 ( .IN1(n3198), .IN2(n5517), .QN(N10479) );
  NAND2X1 U7031 ( .IN1(n5481), .IN2(n5019), .QN(n3199) );
  NOR2X0 U7032 ( .IN1(n3195), .IN2(n5517), .QN(N10480) );
  NAND2X1 U7033 ( .IN1(n5481), .IN2(n5020), .QN(n3196) );
  NOR2X0 U7034 ( .IN1(n3192), .IN2(n5517), .QN(N10481) );
  NAND2X1 U7035 ( .IN1(n5481), .IN2(n5021), .QN(n3193) );
  NOR2X0 U7036 ( .IN1(n3189), .IN2(n5517), .QN(N10482) );
  NAND2X1 U7037 ( .IN1(n5481), .IN2(n5022), .QN(n3190) );
  NOR2X0 U7038 ( .IN1(n3186), .IN2(n5517), .QN(N10483) );
  NAND2X1 U7039 ( .IN1(n5481), .IN2(n5023), .QN(n3187) );
  NOR2X0 U7040 ( .IN1(n3183), .IN2(n5517), .QN(N10484) );
  NAND2X1 U7041 ( .IN1(n5481), .IN2(n5024), .QN(n3184) );
  NOR2X0 U7042 ( .IN1(n2821), .IN2(n5576), .QN(N10605) );
  NAND2X1 U7043 ( .IN1(n5539), .IN2(n4934), .QN(n2822) );
  NOR2X0 U7044 ( .IN1(n2818), .IN2(n5576), .QN(N10606) );
  NAND2X1 U7045 ( .IN1(n5539), .IN2(n4935), .QN(n2819) );
  NOR2X0 U7046 ( .IN1(n2815), .IN2(n5576), .QN(N10607) );
  NAND2X1 U7047 ( .IN1(n5539), .IN2(n4936), .QN(n2816) );
  NOR2X0 U7048 ( .IN1(n2812), .IN2(n5576), .QN(N10608) );
  NAND2X1 U7049 ( .IN1(n5539), .IN2(n4937), .QN(n2813) );
  NOR2X0 U7050 ( .IN1(n2809), .IN2(n5576), .QN(N10609) );
  NAND2X1 U7051 ( .IN1(n5539), .IN2(n4938), .QN(n2810) );
  NOR2X0 U7052 ( .IN1(n2806), .IN2(n5576), .QN(N10610) );
  NAND2X1 U7053 ( .IN1(n5539), .IN2(n4939), .QN(n2807) );
  NOR2X0 U7054 ( .IN1(n2803), .IN2(n5576), .QN(N10611) );
  NAND2X1 U7055 ( .IN1(n5539), .IN2(n4940), .QN(n2804) );
  NOR2X0 U7056 ( .IN1(n2800), .IN2(n5576), .QN(N10612) );
  NAND2X1 U7057 ( .IN1(n5539), .IN2(n4941), .QN(n2801) );
  NOR2X0 U7058 ( .IN1(n2797), .IN2(n5576), .QN(N10613) );
  NAND2X1 U7059 ( .IN1(n5539), .IN2(n4942), .QN(n2798) );
  NOR2X0 U7060 ( .IN1(n2794), .IN2(n5576), .QN(N10614) );
  NAND2X1 U7061 ( .IN1(n5539), .IN2(n4943), .QN(n2795) );
  NOR2X0 U7062 ( .IN1(n2423), .IN2(n5672), .QN(N9684) );
  NAND2X1 U7063 ( .IN1(n5638), .IN2(n5054), .QN(n2424) );
  NOR2X0 U7064 ( .IN1(n2417), .IN2(n5672), .QN(N9685) );
  NAND2X1 U7065 ( .IN1(n5638), .IN2(n5055), .QN(n2418) );
  NOR2X0 U7066 ( .IN1(n2411), .IN2(n5672), .QN(N9686) );
  NAND2X1 U7067 ( .IN1(n5638), .IN2(n5056), .QN(n2412) );
  NOR2X0 U7068 ( .IN1(n2405), .IN2(n5672), .QN(N9687) );
  NAND2X1 U7069 ( .IN1(n5638), .IN2(n5057), .QN(n2406) );
  NOR2X0 U7070 ( .IN1(n2399), .IN2(n5672), .QN(N9688) );
  NAND2X1 U7071 ( .IN1(n5638), .IN2(n5058), .QN(n2400) );
  NOR2X0 U7072 ( .IN1(n2393), .IN2(n5672), .QN(N9689) );
  NAND2X1 U7073 ( .IN1(n5638), .IN2(n5059), .QN(n2394) );
  NOR2X0 U7074 ( .IN1(n2387), .IN2(n5672), .QN(N9690) );
  NAND2X1 U7075 ( .IN1(n5638), .IN2(n5060), .QN(n2388) );
  NOR2X0 U7076 ( .IN1(n2381), .IN2(n5672), .QN(N9691) );
  NAND2X1 U7077 ( .IN1(n5638), .IN2(n5061), .QN(n2382) );
  NOR2X0 U7078 ( .IN1(n2375), .IN2(n5672), .QN(N9692) );
  NAND2X1 U7079 ( .IN1(n5638), .IN2(n5028), .QN(n2376) );
  NOR2X0 U7080 ( .IN1(n2369), .IN2(n5672), .QN(N9693) );
  NAND2X1 U7081 ( .IN1(n5638), .IN2(n5029), .QN(n2370) );
  NOR2X0 U7082 ( .IN1(n2363), .IN2(n5672), .QN(N9694) );
  NAND2X1 U7083 ( .IN1(n5638), .IN2(n5030), .QN(n2364) );
  NOR2X0 U7084 ( .IN1(n2357), .IN2(n5672), .QN(N9695) );
  NAND2X1 U7085 ( .IN1(n5638), .IN2(n5031), .QN(n2358) );
  NOR2X0 U7086 ( .IN1(n1050), .IN2(n5844), .QN(N9943) );
  NAND2X1 U7087 ( .IN1(n5809), .IN2(n5135), .QN(n1051) );
  NOR2X0 U7088 ( .IN1(n1046), .IN2(n5844), .QN(N9944) );
  NAND2X1 U7089 ( .IN1(n5809), .IN2(n5136), .QN(n1047) );
  NOR2X0 U7090 ( .IN1(n1042), .IN2(n5844), .QN(N9945) );
  NAND2X1 U7091 ( .IN1(n5809), .IN2(n5137), .QN(n1043) );
  NOR2X0 U7092 ( .IN1(n1038), .IN2(n5844), .QN(N9946) );
  NAND2X1 U7093 ( .IN1(n5809), .IN2(n5138), .QN(n1039) );
  NOR2X0 U7094 ( .IN1(n1034), .IN2(n5844), .QN(N9947) );
  NAND2X1 U7095 ( .IN1(n5809), .IN2(n5139), .QN(n1035) );
  NOR2X0 U7096 ( .IN1(n1030), .IN2(n5844), .QN(N9948) );
  NAND2X1 U7097 ( .IN1(n5809), .IN2(n5140), .QN(n1031) );
  NOR2X0 U7098 ( .IN1(n1026), .IN2(n5844), .QN(N9949) );
  NAND2X1 U7099 ( .IN1(n5809), .IN2(n5141), .QN(n1027) );
  NOR2X0 U7100 ( .IN1(n1022), .IN2(n5844), .QN(N9950) );
  NAND2X1 U7101 ( .IN1(n5809), .IN2(n5142), .QN(n1023) );
  NOR2X0 U7102 ( .IN1(n1018), .IN2(n5844), .QN(N9951) );
  NAND2X1 U7103 ( .IN1(n5809), .IN2(n5143), .QN(n1019) );
  NOR2X0 U7104 ( .IN1(n1014), .IN2(n5844), .QN(N9952) );
  NAND2X1 U7105 ( .IN1(n5809), .IN2(n5144), .QN(n1015) );
  NOR2X0 U7106 ( .IN1(n1010), .IN2(n5844), .QN(N9953) );
  NAND2X1 U7107 ( .IN1(n5809), .IN2(n5145), .QN(n1011) );
  NOR2X0 U7108 ( .IN1(n1006), .IN2(n5844), .QN(N9954) );
  NAND2X1 U7109 ( .IN1(n5809), .IN2(n5146), .QN(n1007) );
  NOR2X0 U7110 ( .IN1(n4514), .IN2(n5339), .QN(N10073) );
  NAND2X1 U7111 ( .IN1(n5305), .IN2(n5101), .QN(n4515) );
  NOR2X0 U7112 ( .IN1(n4510), .IN2(n5339), .QN(N10074) );
  NAND2X1 U7113 ( .IN1(n5305), .IN2(n5102), .QN(n4511) );
  NOR2X0 U7114 ( .IN1(n4506), .IN2(n5339), .QN(N10075) );
  NAND2X1 U7115 ( .IN1(n5305), .IN2(n5103), .QN(n4507) );
  NOR2X0 U7116 ( .IN1(n4502), .IN2(n5339), .QN(N10076) );
  NAND2X1 U7117 ( .IN1(n5305), .IN2(n5104), .QN(n4503) );
  NOR2X0 U7118 ( .IN1(n4498), .IN2(n5339), .QN(N10077) );
  NAND2X1 U7119 ( .IN1(n5305), .IN2(n5105), .QN(n4499) );
  NOR2X0 U7120 ( .IN1(n4494), .IN2(n5339), .QN(N10078) );
  NAND2X1 U7121 ( .IN1(n5305), .IN2(n5106), .QN(n4495) );
  NOR2X0 U7122 ( .IN1(n4490), .IN2(n5339), .QN(N10079) );
  NAND2X1 U7123 ( .IN1(n5305), .IN2(n5107), .QN(n4491) );
  NOR2X0 U7124 ( .IN1(n4486), .IN2(n5339), .QN(N10080) );
  NAND2X1 U7125 ( .IN1(n5305), .IN2(n5108), .QN(n4487) );
  NOR2X0 U7126 ( .IN1(n4482), .IN2(n5339), .QN(N10081) );
  NAND2X1 U7127 ( .IN1(n5305), .IN2(n5109), .QN(n4483) );
  NOR2X0 U7128 ( .IN1(n4478), .IN2(n5339), .QN(N10082) );
  NAND2X1 U7129 ( .IN1(n5305), .IN2(n5110), .QN(n4479) );
  NOR2X0 U7130 ( .IN1(n4474), .IN2(n5339), .QN(N10083) );
  NAND2X1 U7131 ( .IN1(n5305), .IN2(n5111), .QN(n4475) );
  NOR2X0 U7132 ( .IN1(n4470), .IN2(n5339), .QN(N10084) );
  NAND2X1 U7133 ( .IN1(n5305), .IN2(n5112), .QN(n4471) );
  NOR2X0 U7134 ( .IN1(n4014), .IN2(n5400), .QN(N10203) );
  NAND2X1 U7135 ( .IN1(n5364), .IN2(n4954), .QN(n4015) );
  NOR2X0 U7136 ( .IN1(n4011), .IN2(n5400), .QN(N10204) );
  NAND2X1 U7137 ( .IN1(n5364), .IN2(n4955), .QN(n4012) );
  NOR2X0 U7138 ( .IN1(n4008), .IN2(n5400), .QN(N10205) );
  NAND2X1 U7139 ( .IN1(n5364), .IN2(n4956), .QN(n4009) );
  NOR2X0 U7140 ( .IN1(n4005), .IN2(n5400), .QN(N10206) );
  NAND2X1 U7141 ( .IN1(n5364), .IN2(n4957), .QN(n4006) );
  NOR2X0 U7142 ( .IN1(n4002), .IN2(n5400), .QN(N10207) );
  NAND2X1 U7143 ( .IN1(n5364), .IN2(n4958), .QN(n4003) );
  NOR2X0 U7144 ( .IN1(n3999), .IN2(n5400), .QN(N10208) );
  NAND2X1 U7145 ( .IN1(n5364), .IN2(n4959), .QN(n4000) );
  NOR2X0 U7146 ( .IN1(n3996), .IN2(n5400), .QN(N10209) );
  NAND2X1 U7147 ( .IN1(n5364), .IN2(n4960), .QN(n3997) );
  NOR2X0 U7148 ( .IN1(n3993), .IN2(n5400), .QN(N10210) );
  NAND2X1 U7149 ( .IN1(n5364), .IN2(n4961), .QN(n3994) );
  NOR2X0 U7150 ( .IN1(n3990), .IN2(n5400), .QN(N10211) );
  NAND2X1 U7151 ( .IN1(n5364), .IN2(n4962), .QN(n3991) );
  NOR2X0 U7152 ( .IN1(n3987), .IN2(n5400), .QN(N10212) );
  NAND2X1 U7153 ( .IN1(n5364), .IN2(n4963), .QN(n3988) );
  NOR2X0 U7154 ( .IN1(n3984), .IN2(n5400), .QN(N10213) );
  NAND2X1 U7155 ( .IN1(n5364), .IN2(n5025), .QN(n3985) );
  NOR2X0 U7156 ( .IN1(n3981), .IN2(n5400), .QN(N10214) );
  NAND2X1 U7157 ( .IN1(n5364), .IN2(n4964), .QN(n3982) );
  NOR2X0 U7158 ( .IN1(n3630), .IN2(n5459), .QN(N10333) );
  NAND2X1 U7159 ( .IN1(n5423), .IN2(n4965), .QN(n3631) );
  NOR2X0 U7160 ( .IN1(n3627), .IN2(n5459), .QN(N10334) );
  NAND2X1 U7161 ( .IN1(n5423), .IN2(n4966), .QN(n3628) );
  NOR2X0 U7162 ( .IN1(n3624), .IN2(n5459), .QN(N10335) );
  NAND2X1 U7163 ( .IN1(n5423), .IN2(n4967), .QN(n3625) );
  NOR2X0 U7164 ( .IN1(n3621), .IN2(n5459), .QN(N10336) );
  NAND2X1 U7165 ( .IN1(n5423), .IN2(n4968), .QN(n3622) );
  NOR2X0 U7166 ( .IN1(n3618), .IN2(n5459), .QN(N10337) );
  NAND2X1 U7167 ( .IN1(n5423), .IN2(n4969), .QN(n3619) );
  NOR2X0 U7168 ( .IN1(n3615), .IN2(n5459), .QN(N10338) );
  NAND2X1 U7169 ( .IN1(n5423), .IN2(n4970), .QN(n3616) );
  NOR2X0 U7170 ( .IN1(n3612), .IN2(n5459), .QN(N10339) );
  NAND2X1 U7171 ( .IN1(n5423), .IN2(n4971), .QN(n3613) );
  NOR2X0 U7172 ( .IN1(n3609), .IN2(n5459), .QN(N10340) );
  NAND2X1 U7173 ( .IN1(n5423), .IN2(n4972), .QN(n3610) );
  NOR2X0 U7174 ( .IN1(n3606), .IN2(n5459), .QN(N10341) );
  NAND2X1 U7175 ( .IN1(n5423), .IN2(n4973), .QN(n3607) );
  NOR2X0 U7176 ( .IN1(n3603), .IN2(n5459), .QN(N10342) );
  NAND2X1 U7177 ( .IN1(n5423), .IN2(n4974), .QN(n3604) );
  NOR2X0 U7178 ( .IN1(n3600), .IN2(n5459), .QN(N10343) );
  NAND2X1 U7179 ( .IN1(n5423), .IN2(n5026), .QN(n3601) );
  NOR2X0 U7180 ( .IN1(n3597), .IN2(n5459), .QN(N10344) );
  NAND2X1 U7181 ( .IN1(n5423), .IN2(n4975), .QN(n3598) );
  NOR2X0 U7182 ( .IN1(n3246), .IN2(n5518), .QN(N10463) );
  NAND2X1 U7183 ( .IN1(n5482), .IN2(n4976), .QN(n3247) );
  NOR2X0 U7184 ( .IN1(n3243), .IN2(n5518), .QN(N10464) );
  NAND2X1 U7185 ( .IN1(n5482), .IN2(n4977), .QN(n3244) );
  NOR2X0 U7186 ( .IN1(n3240), .IN2(n5518), .QN(N10465) );
  NAND2X1 U7187 ( .IN1(n5482), .IN2(n4978), .QN(n3241) );
  NOR2X0 U7188 ( .IN1(n3237), .IN2(n5518), .QN(N10466) );
  NAND2X1 U7189 ( .IN1(n5482), .IN2(n4979), .QN(n3238) );
  NOR2X0 U7190 ( .IN1(n3234), .IN2(n5518), .QN(N10467) );
  NAND2X1 U7191 ( .IN1(n5482), .IN2(n4980), .QN(n3235) );
  NOR2X0 U7192 ( .IN1(n3231), .IN2(n5518), .QN(N10468) );
  NAND2X1 U7193 ( .IN1(n5482), .IN2(n4981), .QN(n3232) );
  NOR2X0 U7194 ( .IN1(n3228), .IN2(n5518), .QN(N10469) );
  NAND2X1 U7195 ( .IN1(n5482), .IN2(n4982), .QN(n3229) );
  NOR2X0 U7196 ( .IN1(n3225), .IN2(n5518), .QN(N10470) );
  NAND2X1 U7197 ( .IN1(n5482), .IN2(n4983), .QN(n3226) );
  NOR2X0 U7198 ( .IN1(n3222), .IN2(n5518), .QN(N10471) );
  NAND2X1 U7199 ( .IN1(n5482), .IN2(n4984), .QN(n3223) );
  NOR2X0 U7200 ( .IN1(n3219), .IN2(n5518), .QN(N10472) );
  NAND2X1 U7201 ( .IN1(n5482), .IN2(n4985), .QN(n3220) );
  NOR2X0 U7202 ( .IN1(n3216), .IN2(n5518), .QN(N10473) );
  NAND2X1 U7203 ( .IN1(n5482), .IN2(n5027), .QN(n3217) );
  NOR2X0 U7204 ( .IN1(n3213), .IN2(n5518), .QN(N10474) );
  NAND2X1 U7205 ( .IN1(n5482), .IN2(n4986), .QN(n3214) );
  NOR2X0 U7206 ( .IN1(n2857), .IN2(n5577), .QN(N10593) );
  NAND2X1 U7207 ( .IN1(n5540), .IN2(n4923), .QN(n2858) );
  NOR2X0 U7208 ( .IN1(n2854), .IN2(n5577), .QN(N10594) );
  NAND2X1 U7209 ( .IN1(n5540), .IN2(n4924), .QN(n2855) );
  NOR2X0 U7210 ( .IN1(n2851), .IN2(n5577), .QN(N10595) );
  NAND2X1 U7211 ( .IN1(n5540), .IN2(n4925), .QN(n2852) );
  NOR2X0 U7212 ( .IN1(n2848), .IN2(n5577), .QN(N10596) );
  NAND2X1 U7213 ( .IN1(n5540), .IN2(n4926), .QN(n2849) );
  NOR2X0 U7214 ( .IN1(n2845), .IN2(n5577), .QN(N10597) );
  NAND2X1 U7215 ( .IN1(n5540), .IN2(n4927), .QN(n2846) );
  NOR2X0 U7216 ( .IN1(n2842), .IN2(n5577), .QN(N10598) );
  NAND2X1 U7217 ( .IN1(n5540), .IN2(n4928), .QN(n2843) );
  NOR2X0 U7218 ( .IN1(n2839), .IN2(n5577), .QN(N10599) );
  NAND2X1 U7219 ( .IN1(n5540), .IN2(n4929), .QN(n2840) );
  NOR2X0 U7220 ( .IN1(n2836), .IN2(n5577), .QN(N10600) );
  NAND2X1 U7221 ( .IN1(n5540), .IN2(n4987), .QN(n2837) );
  NOR2X0 U7222 ( .IN1(n2833), .IN2(n5577), .QN(N10601) );
  NAND2X1 U7223 ( .IN1(n5540), .IN2(n4930), .QN(n2834) );
  NOR2X0 U7224 ( .IN1(n2830), .IN2(n5577), .QN(N10602) );
  NAND2X1 U7225 ( .IN1(n5540), .IN2(n4931), .QN(n2831) );
  NOR2X0 U7226 ( .IN1(n2827), .IN2(n5577), .QN(N10603) );
  NAND2X1 U7227 ( .IN1(n5540), .IN2(n4944), .QN(n2828) );
  NOR2X0 U7228 ( .IN1(n2824), .IN2(n5577), .QN(N10604) );
  NAND2X1 U7229 ( .IN1(n5540), .IN2(n4932), .QN(n2825) );
  NOR2X0 U7230 ( .IN1(n2351), .IN2(n5671), .QN(N9696) );
  NAND2X1 U7231 ( .IN1(n5637), .IN2(n5032), .QN(n2352) );
  NOR2X0 U7232 ( .IN1(n2345), .IN2(n5671), .QN(N9697) );
  NAND2X1 U7233 ( .IN1(n5637), .IN2(n5033), .QN(n2346) );
  NOR2X0 U7234 ( .IN1(n2339), .IN2(n5671), .QN(N9698) );
  NAND2X1 U7235 ( .IN1(n5637), .IN2(n5034), .QN(n2340) );
  NOR2X0 U7236 ( .IN1(n2333), .IN2(n5671), .QN(N9699) );
  NAND2X1 U7237 ( .IN1(n5637), .IN2(n5035), .QN(n2334) );
  NOR2X0 U7238 ( .IN1(n2327), .IN2(n5671), .QN(N9700) );
  NAND2X1 U7239 ( .IN1(n5637), .IN2(n5036), .QN(n2328) );
  NOR2X0 U7240 ( .IN1(n2321), .IN2(n5671), .QN(N9701) );
  NAND2X1 U7241 ( .IN1(n5637), .IN2(n5037), .QN(n2322) );
  NOR2X0 U7242 ( .IN1(n2315), .IN2(n5671), .QN(N9702) );
  NAND2X1 U7243 ( .IN1(n5637), .IN2(n5038), .QN(n2316) );
  NOR2X0 U7244 ( .IN1(n2309), .IN2(n5671), .QN(N9703) );
  NAND2X1 U7245 ( .IN1(n5637), .IN2(n5039), .QN(n2310) );
  NOR2X0 U7246 ( .IN1(n2303), .IN2(n5671), .QN(N9704) );
  NAND2X1 U7247 ( .IN1(n5637), .IN2(n5040), .QN(n2304) );
  NOR2X0 U7248 ( .IN1(n2297), .IN2(n5671), .QN(N9705) );
  NAND2X1 U7249 ( .IN1(n5637), .IN2(n5041), .QN(n2298) );
  NOR2X0 U7250 ( .IN1(n4466), .IN2(n5338), .QN(N10085) );
  NAND2X1 U7251 ( .IN1(n5304), .IN2(n5113), .QN(n4467) );
  NOR2X0 U7252 ( .IN1(n4462), .IN2(n5338), .QN(N10086) );
  NAND2X1 U7253 ( .IN1(n5304), .IN2(n5114), .QN(n4463) );
  NOR2X0 U7254 ( .IN1(n4458), .IN2(n5338), .QN(N10087) );
  NAND2X1 U7255 ( .IN1(n5304), .IN2(n5115), .QN(n4459) );
  NOR2X0 U7256 ( .IN1(n4454), .IN2(n5338), .QN(N10088) );
  NAND2X1 U7257 ( .IN1(n5304), .IN2(n5116), .QN(n4455) );
  NOR2X0 U7258 ( .IN1(n4450), .IN2(n5338), .QN(N10089) );
  NAND2X1 U7259 ( .IN1(n5304), .IN2(n5117), .QN(n4451) );
  NOR2X0 U7260 ( .IN1(n4446), .IN2(n5338), .QN(N10090) );
  NAND2X1 U7261 ( .IN1(n5304), .IN2(n5118), .QN(n4447) );
  NOR2X0 U7262 ( .IN1(n4442), .IN2(n5338), .QN(N10091) );
  NAND2X1 U7263 ( .IN1(n5304), .IN2(n5119), .QN(n4443) );
  NOR2X0 U7264 ( .IN1(n4438), .IN2(n5338), .QN(N10092) );
  NAND2X1 U7265 ( .IN1(n5304), .IN2(n5120), .QN(n4439) );
  NOR2X0 U7266 ( .IN1(n4434), .IN2(n5338), .QN(N10093) );
  NAND2X1 U7267 ( .IN1(n5304), .IN2(n5121), .QN(n4435) );
  NOR2X0 U7268 ( .IN1(n4430), .IN2(n5338), .QN(N10094) );
  NAND2X1 U7269 ( .IN1(n5304), .IN2(n5122), .QN(n4431) );
  NOR2X0 U7270 ( .IN1(n1002), .IN2(n5843), .QN(N9955) );
  NAND2X1 U7271 ( .IN1(n5808), .IN2(n5147), .QN(n1003) );
  NOR2X0 U7272 ( .IN1(n998), .IN2(n5843), .QN(N9956) );
  NAND2X1 U7273 ( .IN1(n5808), .IN2(n5148), .QN(n999) );
  NOR2X0 U7274 ( .IN1(n994), .IN2(n5843), .QN(N9957) );
  NAND2X1 U7275 ( .IN1(n5808), .IN2(n5149), .QN(n995) );
  NOR2X0 U7276 ( .IN1(n990), .IN2(n5843), .QN(N9958) );
  NAND2X1 U7277 ( .IN1(n5808), .IN2(n5150), .QN(n991) );
  NOR2X0 U7278 ( .IN1(n986), .IN2(n5843), .QN(N9959) );
  NAND2X1 U7279 ( .IN1(n5808), .IN2(n5151), .QN(n987) );
  NOR2X0 U7280 ( .IN1(n982), .IN2(n5843), .QN(N9960) );
  NAND2X1 U7281 ( .IN1(n5808), .IN2(n5152), .QN(n983) );
  NOR2X0 U7282 ( .IN1(n978), .IN2(n5843), .QN(N9961) );
  NAND2X1 U7283 ( .IN1(n5808), .IN2(n5153), .QN(n979) );
  NOR2X0 U7284 ( .IN1(n974), .IN2(n5843), .QN(N9962) );
  NAND2X1 U7285 ( .IN1(n5808), .IN2(n5154), .QN(n975) );
  NOR2X0 U7286 ( .IN1(n970), .IN2(n5843), .QN(N9963) );
  NAND2X1 U7287 ( .IN1(n5808), .IN2(n5155), .QN(n971) );
  NOR2X0 U7288 ( .IN1(n966), .IN2(n5843), .QN(N9964) );
  NAND2X1 U7289 ( .IN1(n5808), .IN2(n5156), .QN(n967) );
  INVX0 U7290 ( .INP(\decodedPacket[4][107] ), .ZN(n6208) );
  INVX0 U7291 ( .INP(\decodedPacket[4][108] ), .ZN(n6209) );
  INVX0 U7292 ( .INP(\decodedPacket[4][109] ), .ZN(n6210) );
  INVX0 U7293 ( .INP(\decodedPacket[4][110] ), .ZN(n6211) );
  INVX0 U7294 ( .INP(\decodedPacket[4][111] ), .ZN(n6212) );
  INVX0 U7295 ( .INP(\decodedPacket[6][107] ), .ZN(n6362) );
  INVX0 U7296 ( .INP(\decodedPacket[6][108] ), .ZN(n6363) );
  INVX0 U7297 ( .INP(\decodedPacket[6][109] ), .ZN(n6364) );
  INVX0 U7298 ( .INP(\decodedPacket[6][110] ), .ZN(n6365) );
  INVX0 U7299 ( .INP(\decodedPacket[6][111] ), .ZN(n6366) );
  INVX0 U7300 ( .INP(\decodedPacket[4][85] ), .ZN(n6200) );
  INVX0 U7301 ( .INP(\decodedPacket[4][86] ), .ZN(n6201) );
  INVX0 U7302 ( .INP(\decodedPacket[4][87] ), .ZN(n6202) );
  INVX0 U7303 ( .INP(\decodedPacket[4][88] ), .ZN(n6203) );
  INVX0 U7304 ( .INP(\decodedPacket[4][89] ), .ZN(n6204) );
  INVX0 U7305 ( .INP(\decodedPacket[4][90] ), .ZN(n6205) );
  INVX0 U7306 ( .INP(\decodedPacket[6][85] ), .ZN(n6354) );
  INVX0 U7307 ( .INP(\decodedPacket[6][86] ), .ZN(n6355) );
  INVX0 U7308 ( .INP(\decodedPacket[6][87] ), .ZN(n6356) );
  INVX0 U7309 ( .INP(\decodedPacket[6][88] ), .ZN(n6357) );
  INVX0 U7310 ( .INP(\decodedPacket[6][89] ), .ZN(n6358) );
  INVX0 U7311 ( .INP(\decodedPacket[6][90] ), .ZN(n6359) );
  INVX0 U7312 ( .INP(\decodedPacket[4][73] ), .ZN(n6251) );
  INVX0 U7313 ( .INP(\decodedPacket[4][74] ), .ZN(n6250) );
  INVX0 U7314 ( .INP(\decodedPacket[4][75] ), .ZN(n6249) );
  INVX0 U7315 ( .INP(\decodedPacket[4][76] ), .ZN(n6248) );
  INVX0 U7316 ( .INP(\decodedPacket[6][73] ), .ZN(n6405) );
  INVX0 U7317 ( .INP(\decodedPacket[6][74] ), .ZN(n6404) );
  INVX0 U7318 ( .INP(\decodedPacket[6][75] ), .ZN(n6403) );
  INVX0 U7319 ( .INP(\decodedPacket[6][76] ), .ZN(n6402) );
  INVX0 U7320 ( .INP(\decodedPacket[4][83] ), .ZN(n6261) );
  INVX0 U7321 ( .INP(\decodedPacket[4][94] ), .ZN(n6265) );
  INVX0 U7322 ( .INP(\decodedPacket[4][95] ), .ZN(n6266) );
  INVX0 U7323 ( .INP(\decodedPacket[6][83] ), .ZN(n6415) );
  INVX0 U7324 ( .INP(\decodedPacket[6][94] ), .ZN(n6419) );
  INVX0 U7325 ( .INP(\decodedPacket[6][95] ), .ZN(n6420) );
  INVX0 U7326 ( .INP(\decodedPacket[4][92] ), .ZN(n6263) );
  INVX0 U7327 ( .INP(\decodedPacket[4][96] ), .ZN(n6267) );
  INVX0 U7328 ( .INP(\decodedPacket[6][92] ), .ZN(n6417) );
  INVX0 U7329 ( .INP(\decodedPacket[6][96] ), .ZN(n6421) );
  INVX0 U7330 ( .INP(\decodedPacket[4][78] ), .ZN(n6256) );
  INVX0 U7331 ( .INP(\decodedPacket[4][93] ), .ZN(n6264) );
  INVX0 U7332 ( .INP(\decodedPacket[6][78] ), .ZN(n6410) );
  INVX0 U7333 ( .INP(\decodedPacket[6][93] ), .ZN(n6418) );
  INVX0 U7334 ( .INP(\decodedPacket[3][78] ), .ZN(n6093) );
  INVX0 U7335 ( .INP(\decodedPacket[3][83] ), .ZN(n6092) );
  INVX0 U7336 ( .INP(\decodedPacket[4][71] ), .ZN(n6206) );
  INVX0 U7337 ( .INP(\decodedPacket[6][71] ), .ZN(n6360) );
  INVX0 U7338 ( .INP(\decodedPacket[5][78] ), .ZN(n6247) );
  INVX0 U7339 ( .INP(\decodedPacket[5][83] ), .ZN(n6246) );
  INVX0 U7340 ( .INP(\decodedPacket[3][92] ), .ZN(n6074) );
  INVX0 U7341 ( .INP(\decodedPacket[3][97] ), .ZN(n6069) );
  INVX0 U7342 ( .INP(\decodedPacket[5][92] ), .ZN(n6228) );
  INVX0 U7343 ( .INP(\decodedPacket[5][97] ), .ZN(n6223) );
  INVX0 U7344 ( .INP(\decodedPacket[3][93] ), .ZN(n6073) );
  INVX0 U7345 ( .INP(\decodedPacket[3][94] ), .ZN(n6072) );
  INVX0 U7346 ( .INP(\decodedPacket[3][95] ), .ZN(n6071) );
  INVX0 U7347 ( .INP(\decodedPacket[3][96] ), .ZN(n6070) );
  INVX0 U7348 ( .INP(\decodedPacket[5][93] ), .ZN(n6227) );
  INVX0 U7349 ( .INP(\decodedPacket[5][94] ), .ZN(n6226) );
  INVX0 U7350 ( .INP(\decodedPacket[5][95] ), .ZN(n6225) );
  INVX0 U7351 ( .INP(\decodedPacket[5][96] ), .ZN(n6224) );
  INVX0 U7352 ( .INP(\decodedPacket[7][78] ), .ZN(n6401) );
  INVX0 U7353 ( .INP(\decodedPacket[7][83] ), .ZN(n6400) );
  INVX0 U7354 ( .INP(\decodedPacket[7][92] ), .ZN(n6382) );
  INVX0 U7355 ( .INP(\decodedPacket[7][97] ), .ZN(n6377) );
  INVX0 U7356 ( .INP(\decodedPacket[7][93] ), .ZN(n6381) );
  INVX0 U7357 ( .INP(\decodedPacket[7][94] ), .ZN(n6380) );
  INVX0 U7358 ( .INP(\decodedPacket[7][95] ), .ZN(n6379) );
  INVX0 U7359 ( .INP(\decodedPacket[7][96] ), .ZN(n6378) );
  OAI22X1 U7360 ( .IN1(n5606), .IN2(n2380), .IN3(n6025), .IN4(n5608), .QN(
        n5202) );
  OAI22X1 U7361 ( .IN1(n5606), .IN2(n2374), .IN3(n6024), .IN4(n5614), .QN(
        n5203) );
  OAI22X1 U7362 ( .IN1(n5606), .IN2(n2368), .IN3(n6023), .IN4(n5597), .QN(
        n5204) );
  OAI22X1 U7363 ( .IN1(n5606), .IN2(n2362), .IN3(n6022), .IN4(n5609), .QN(
        n5205) );
  OAI22X1 U7364 ( .IN1(n5606), .IN2(n2356), .IN3(n6021), .IN4(n5612), .QN(
        n5206) );
  OAI22X1 U7365 ( .IN1(n5606), .IN2(n2350), .IN3(n6020), .IN4(n5597), .QN(
        n5207) );
  OAI22X1 U7366 ( .IN1(n5606), .IN2(n2344), .IN3(n6019), .IN4(n5598), .QN(
        n5208) );
  OAI22X1 U7367 ( .IN1(n5606), .IN2(n2338), .IN3(n6018), .IN4(n5599), .QN(
        n5209) );
  OAI22X1 U7368 ( .IN1(n5606), .IN2(n2332), .IN3(n6017), .IN4(n5610), .QN(
        n5210) );
  OAI22X1 U7369 ( .IN1(n5606), .IN2(n2326), .IN3(n6016), .IN4(n5613), .QN(
        n5211) );
  OAI22X1 U7370 ( .IN1(n5605), .IN2(n2320), .IN3(n6015), .IN4(n5614), .QN(
        n5212) );
  OAI22X1 U7371 ( .IN1(n5605), .IN2(n2314), .IN3(n6014), .IN4(n5615), .QN(
        n5213) );
  OAI22X1 U7372 ( .IN1(n5605), .IN2(n2308), .IN3(n6013), .IN4(n5613), .QN(
        n5214) );
  OAI22X1 U7373 ( .IN1(n5605), .IN2(n2302), .IN3(n6012), .IN4(n5597), .QN(
        n5215) );
  INVX0 U7374 ( .INP(\decodedPacket[2][12] ), .ZN(n6036) );
  INVX0 U7375 ( .INP(\decodedPacket[2][13] ), .ZN(n6035) );
  INVX0 U7376 ( .INP(\decodedPacket[2][14] ), .ZN(n6034) );
  INVX0 U7377 ( .INP(\decodedPacket[2][15] ), .ZN(n6033) );
  INVX0 U7378 ( .INP(\decodedPacket[2][16] ), .ZN(n6032) );
  INVX0 U7379 ( .INP(\decodedPacket[2][5] ), .ZN(n6011) );
  INVX0 U7380 ( .INP(\decodedPacket[2][6] ), .ZN(n6010) );
  INVX0 U7381 ( .INP(\decodedPacket[2][7] ), .ZN(n6009) );
  INVX0 U7382 ( .INP(\decodedPacket[2][8] ), .ZN(n6008) );
  INVX0 U7383 ( .INP(\decodedPacket[2][9] ), .ZN(n6007) );
  INVX0 U7384 ( .INP(\decodedPacket[2][11] ), .ZN(n6037) );
  INVX0 U7385 ( .INP(\decodedPacket[2][30] ), .ZN(n6018) );
  INVX0 U7386 ( .INP(\decodedPacket[2][10] ), .ZN(n6038) );
  INVX0 U7387 ( .INP(\decodedPacket[2][17] ), .ZN(n6031) );
  INVX0 U7388 ( .INP(\decodedPacket[2][18] ), .ZN(n6030) );
  INVX0 U7389 ( .INP(\decodedPacket[2][19] ), .ZN(n6029) );
  INVX0 U7390 ( .INP(\decodedPacket[2][20] ), .ZN(n6028) );
  INVX0 U7391 ( .INP(\decodedPacket[2][21] ), .ZN(n6027) );
  INVX0 U7392 ( .INP(\decodedPacket[2][22] ), .ZN(n6026) );
  INVX0 U7393 ( .INP(\decodedPacket[2][23] ), .ZN(n6025) );
  INVX0 U7394 ( .INP(\decodedPacket[2][24] ), .ZN(n6024) );
  INVX0 U7395 ( .INP(\decodedPacket[2][25] ), .ZN(n6023) );
  INVX0 U7396 ( .INP(\decodedPacket[2][26] ), .ZN(n6022) );
  INVX0 U7397 ( .INP(\decodedPacket[2][27] ), .ZN(n6021) );
  INVX0 U7398 ( .INP(\decodedPacket[2][28] ), .ZN(n6020) );
  INVX0 U7399 ( .INP(\decodedPacket[2][29] ), .ZN(n6019) );
  OAI22X1 U7400 ( .IN1(n5607), .IN2(n2488), .IN3(n6011), .IN4(n5599), .QN(
        n5216) );
  OAI22X1 U7401 ( .IN1(n5607), .IN2(n2482), .IN3(n6010), .IN4(n5614), .QN(
        n5217) );
  OAI22X1 U7402 ( .IN1(n5607), .IN2(n2476), .IN3(n6009), .IN4(n5611), .QN(
        n5218) );
  OAI22X1 U7403 ( .IN1(n5607), .IN2(n2470), .IN3(n6008), .IN4(n5612), .QN(
        n5219) );
  OAI22X1 U7404 ( .IN1(n5607), .IN2(n2464), .IN3(n6007), .IN4(n5597), .QN(
        n5220) );
  OAI22X1 U7405 ( .IN1(n5607), .IN2(n2458), .IN3(n6038), .IN4(n5614), .QN(
        n5221) );
  OAI22X1 U7406 ( .IN1(n5607), .IN2(n2452), .IN3(n6037), .IN4(n5615), .QN(
        n5222) );
  OAI22X1 U7407 ( .IN1(n5607), .IN2(n2446), .IN3(n6036), .IN4(n5608), .QN(
        n5223) );
  OAI22X1 U7408 ( .IN1(n5607), .IN2(n2440), .IN3(n6035), .IN4(n5608), .QN(
        n5224) );
  OAI22X1 U7409 ( .IN1(n5607), .IN2(n2434), .IN3(n6034), .IN4(n5609), .QN(
        n5225) );
  OAI22X1 U7410 ( .IN1(n5607), .IN2(n2428), .IN3(n6033), .IN4(n5610), .QN(
        n5226) );
  OAI22X1 U7411 ( .IN1(n5607), .IN2(n2422), .IN3(n6032), .IN4(n5614), .QN(
        n5227) );
  OAI22X1 U7412 ( .IN1(n5607), .IN2(n2416), .IN3(n6031), .IN4(n5613), .QN(
        n5228) );
  OAI22X1 U7413 ( .IN1(n5606), .IN2(n2410), .IN3(n6030), .IN4(n5615), .QN(
        n5229) );
  OAI22X1 U7414 ( .IN1(n5606), .IN2(n2404), .IN3(n6029), .IN4(n5611), .QN(
        n5230) );
  OAI22X1 U7415 ( .IN1(n5606), .IN2(n2398), .IN3(n6028), .IN4(n5599), .QN(
        n5231) );
  OAI22X1 U7416 ( .IN1(n5606), .IN2(n2392), .IN3(n6027), .IN4(n5613), .QN(
        n5232) );
  OAI22X1 U7417 ( .IN1(n5606), .IN2(n2386), .IN3(n6026), .IN4(n5611), .QN(
        n5233) );
  INVX0 U7418 ( .INP(\decodedPacket[2][31] ), .ZN(n6017) );
  INVX0 U7419 ( .INP(\decodedPacket[2][32] ), .ZN(n6016) );
  INVX0 U7420 ( .INP(\decodedPacket[2][33] ), .ZN(n6015) );
  INVX0 U7421 ( .INP(\decodedPacket[2][34] ), .ZN(n6014) );
  INVX0 U7422 ( .INP(\decodedPacket[2][35] ), .ZN(n6013) );
  INVX0 U7423 ( .INP(\decodedPacket[2][36] ), .ZN(n6012) );
  INVX0 U7424 ( .INP(\decodedPacket[2][112] ), .ZN(n6059) );
  INVX0 U7425 ( .INP(\decodedPacket[2][113] ), .ZN(n6060) );
  INVX0 U7426 ( .INP(\decodedPacket[2][114] ), .ZN(n6061) );
  NAND2X1 U7427 ( .IN1(n5775), .IN2(\decodedPacket[2][5] ), .QN(n1093) );
  NAND2X1 U7428 ( .IN1(n5775), .IN2(\decodedPacket[2][6] ), .QN(n1089) );
  NAND2X1 U7429 ( .IN1(n5775), .IN2(\decodedPacket[2][7] ), .QN(n1085) );
  NAND2X1 U7430 ( .IN1(n5775), .IN2(\decodedPacket[2][8] ), .QN(n1081) );
  NAND2X1 U7431 ( .IN1(n5775), .IN2(\decodedPacket[2][9] ), .QN(n1077) );
  NAND2X1 U7432 ( .IN1(n5775), .IN2(\decodedPacket[2][10] ), .QN(n1073) );
  NAND2X1 U7433 ( .IN1(n5775), .IN2(\decodedPacket[2][11] ), .QN(n1069) );
  NAND2X1 U7434 ( .IN1(n5775), .IN2(\decodedPacket[2][12] ), .QN(n1065) );
  NAND2X1 U7435 ( .IN1(n5775), .IN2(\decodedPacket[2][13] ), .QN(n1061) );
  NAND2X1 U7436 ( .IN1(n5775), .IN2(\decodedPacket[2][14] ), .QN(n1057) );
  NAND2X1 U7437 ( .IN1(n5774), .IN2(\decodedPacket[2][15] ), .QN(n1053) );
  NAND2X1 U7438 ( .IN1(n5774), .IN2(\decodedPacket[2][16] ), .QN(n1049) );
  NAND2X1 U7439 ( .IN1(n5774), .IN2(\decodedPacket[2][17] ), .QN(n1045) );
  NAND2X1 U7440 ( .IN1(n5774), .IN2(\decodedPacket[2][18] ), .QN(n1041) );
  NAND2X1 U7441 ( .IN1(n5774), .IN2(\decodedPacket[2][19] ), .QN(n1037) );
  NAND2X1 U7442 ( .IN1(n5774), .IN2(\decodedPacket[2][20] ), .QN(n1033) );
  NAND2X1 U7443 ( .IN1(n5774), .IN2(\decodedPacket[2][21] ), .QN(n1029) );
  NAND2X1 U7444 ( .IN1(n5774), .IN2(\decodedPacket[2][22] ), .QN(n1025) );
  NAND2X1 U7445 ( .IN1(n5774), .IN2(\decodedPacket[2][23] ), .QN(n1021) );
  NAND2X1 U7446 ( .IN1(n5774), .IN2(\decodedPacket[2][24] ), .QN(n1017) );
  NAND2X1 U7447 ( .IN1(n5774), .IN2(\decodedPacket[2][25] ), .QN(n1013) );
  NAND2X1 U7448 ( .IN1(n5774), .IN2(\decodedPacket[2][26] ), .QN(n1009) );
  NAND2X1 U7449 ( .IN1(n5773), .IN2(\decodedPacket[2][27] ), .QN(n1005) );
  NAND2X1 U7450 ( .IN1(n5773), .IN2(\decodedPacket[2][28] ), .QN(n1001) );
  NAND2X1 U7451 ( .IN1(n5773), .IN2(\decodedPacket[2][29] ), .QN(n997) );
  NAND2X1 U7452 ( .IN1(n5773), .IN2(\decodedPacket[2][30] ), .QN(n993) );
  NAND2X1 U7453 ( .IN1(n5773), .IN2(\decodedPacket[2][31] ), .QN(n989) );
  NAND2X1 U7454 ( .IN1(n5773), .IN2(\decodedPacket[2][32] ), .QN(n985) );
  NAND2X1 U7455 ( .IN1(n5773), .IN2(\decodedPacket[2][33] ), .QN(n981) );
  NAND2X1 U7456 ( .IN1(n5773), .IN2(\decodedPacket[2][34] ), .QN(n977) );
  NAND2X1 U7457 ( .IN1(n5773), .IN2(\decodedPacket[2][35] ), .QN(n973) );
  NAND2X1 U7458 ( .IN1(n5773), .IN2(\decodedPacket[2][36] ), .QN(n969) );
  NAND2X1 U7459 ( .IN1(n5278), .IN2(\decodedPacket[2][5] ), .QN(n4557) );
  NAND2X1 U7460 ( .IN1(n5278), .IN2(\decodedPacket[2][6] ), .QN(n4553) );
  NAND2X1 U7461 ( .IN1(n5278), .IN2(\decodedPacket[2][7] ), .QN(n4549) );
  NAND2X1 U7462 ( .IN1(n5278), .IN2(\decodedPacket[2][8] ), .QN(n4545) );
  NAND2X1 U7463 ( .IN1(n5278), .IN2(\decodedPacket[2][9] ), .QN(n4541) );
  NAND2X1 U7464 ( .IN1(n5278), .IN2(\decodedPacket[2][10] ), .QN(n4537) );
  NAND2X1 U7465 ( .IN1(n5278), .IN2(\decodedPacket[2][11] ), .QN(n4533) );
  NAND2X1 U7466 ( .IN1(n5278), .IN2(\decodedPacket[2][12] ), .QN(n4529) );
  NAND2X1 U7467 ( .IN1(n5278), .IN2(\decodedPacket[2][13] ), .QN(n4525) );
  NAND2X1 U7468 ( .IN1(n5278), .IN2(\decodedPacket[2][14] ), .QN(n4521) );
  NAND2X1 U7469 ( .IN1(n5277), .IN2(\decodedPacket[2][15] ), .QN(n4517) );
  NAND2X1 U7470 ( .IN1(n5277), .IN2(\decodedPacket[2][16] ), .QN(n4513) );
  NAND2X1 U7471 ( .IN1(n5277), .IN2(\decodedPacket[2][17] ), .QN(n4509) );
  NAND2X1 U7472 ( .IN1(n5277), .IN2(\decodedPacket[2][18] ), .QN(n4505) );
  NAND2X1 U7473 ( .IN1(n5277), .IN2(\decodedPacket[2][19] ), .QN(n4501) );
  NAND2X1 U7474 ( .IN1(n5277), .IN2(\decodedPacket[2][20] ), .QN(n4497) );
  NAND2X1 U7475 ( .IN1(n5277), .IN2(\decodedPacket[2][21] ), .QN(n4493) );
  NAND2X1 U7476 ( .IN1(n5277), .IN2(\decodedPacket[2][22] ), .QN(n4489) );
  NAND2X1 U7477 ( .IN1(n5277), .IN2(\decodedPacket[2][23] ), .QN(n4485) );
  NAND2X1 U7478 ( .IN1(n5277), .IN2(\decodedPacket[2][24] ), .QN(n4481) );
  NAND2X1 U7479 ( .IN1(n5277), .IN2(\decodedPacket[2][25] ), .QN(n4477) );
  NAND2X1 U7480 ( .IN1(n5277), .IN2(\decodedPacket[2][26] ), .QN(n4473) );
  NAND2X1 U7481 ( .IN1(n5276), .IN2(\decodedPacket[2][27] ), .QN(n4469) );
  NAND2X1 U7482 ( .IN1(n5276), .IN2(\decodedPacket[2][28] ), .QN(n4465) );
  NAND2X1 U7483 ( .IN1(n5276), .IN2(\decodedPacket[2][29] ), .QN(n4461) );
  NAND2X1 U7484 ( .IN1(n5276), .IN2(\decodedPacket[2][30] ), .QN(n4457) );
  NAND2X1 U7485 ( .IN1(n5276), .IN2(\decodedPacket[2][31] ), .QN(n4453) );
  NAND2X1 U7486 ( .IN1(n5276), .IN2(\decodedPacket[2][32] ), .QN(n4449) );
  NAND2X1 U7487 ( .IN1(n5276), .IN2(\decodedPacket[2][33] ), .QN(n4445) );
  NAND2X1 U7488 ( .IN1(n5276), .IN2(\decodedPacket[2][34] ), .QN(n4441) );
  NAND2X1 U7489 ( .IN1(n5276), .IN2(\decodedPacket[2][35] ), .QN(n4437) );
  NAND2X1 U7490 ( .IN1(n5276), .IN2(\decodedPacket[2][36] ), .QN(n4433) );
  AND2X1 U7491 ( .IN1(\decodedPacket[2][12] ), .IN2(n5693), .Q(n5234) );
  AND2X1 U7492 ( .IN1(\decodedPacket[2][13] ), .IN2(n5693), .Q(n5235) );
  AND2X1 U7493 ( .IN1(\decodedPacket[2][14] ), .IN2(n5693), .Q(n5236) );
  AND2X1 U7494 ( .IN1(\decodedPacket[2][15] ), .IN2(n5692), .Q(n5237) );
  AND2X1 U7495 ( .IN1(\decodedPacket[2][16] ), .IN2(n5692), .Q(n5238) );
  AND2X1 U7496 ( .IN1(\decodedPacket[2][17] ), .IN2(n5692), .Q(n5239) );
  AND2X1 U7497 ( .IN1(\decodedPacket[2][18] ), .IN2(n5692), .Q(n5240) );
  AND2X1 U7498 ( .IN1(\decodedPacket[2][19] ), .IN2(n5692), .Q(n5241) );
  AND2X1 U7499 ( .IN1(\decodedPacket[2][20] ), .IN2(n5692), .Q(n5242) );
  AND2X1 U7500 ( .IN1(\decodedPacket[2][21] ), .IN2(n5692), .Q(n5243) );
  AND2X1 U7501 ( .IN1(\decodedPacket[2][22] ), .IN2(n5692), .Q(n5244) );
  AND2X1 U7502 ( .IN1(\decodedPacket[2][23] ), .IN2(n5692), .Q(n5245) );
  AND2X1 U7503 ( .IN1(\decodedPacket[2][24] ), .IN2(n5692), .Q(n5246) );
  AND2X1 U7504 ( .IN1(\decodedPacket[2][25] ), .IN2(n5692), .Q(n5247) );
  AND2X1 U7505 ( .IN1(\decodedPacket[2][26] ), .IN2(n5692), .Q(n5248) );
  AND2X1 U7506 ( .IN1(\decodedPacket[2][27] ), .IN2(n5691), .Q(n5249) );
  AND2X1 U7507 ( .IN1(\decodedPacket[2][28] ), .IN2(n5691), .Q(n5250) );
  AND2X1 U7508 ( .IN1(\decodedPacket[2][29] ), .IN2(n5691), .Q(n5251) );
  AND2X1 U7509 ( .IN1(\decodedPacket[2][30] ), .IN2(n5691), .Q(n5252) );
  AND2X1 U7510 ( .IN1(\decodedPacket[2][31] ), .IN2(n5691), .Q(n5253) );
  AND2X1 U7511 ( .IN1(\decodedPacket[2][32] ), .IN2(n5691), .Q(n5254) );
  AND2X1 U7512 ( .IN1(\decodedPacket[2][33] ), .IN2(n5691), .Q(n5255) );
  AND2X1 U7513 ( .IN1(\decodedPacket[2][34] ), .IN2(n5691), .Q(n5256) );
  AND2X1 U7514 ( .IN1(\decodedPacket[2][35] ), .IN2(n5691), .Q(n5257) );
  AND2X1 U7515 ( .IN1(\decodedPacket[2][36] ), .IN2(n5691), .Q(n5258) );
  AND2X1 U7516 ( .IN1(\decodedPacket[2][5] ), .IN2(n5693), .Q(n5259) );
  AND2X1 U7517 ( .IN1(\decodedPacket[2][6] ), .IN2(n5693), .Q(n5260) );
  AND2X1 U7518 ( .IN1(\decodedPacket[2][7] ), .IN2(n5693), .Q(n5261) );
  AND2X1 U7519 ( .IN1(\decodedPacket[2][8] ), .IN2(n5693), .Q(n5262) );
  AND2X1 U7520 ( .IN1(\decodedPacket[2][9] ), .IN2(n5693), .Q(n5263) );
  AND2X1 U7521 ( .IN1(\decodedPacket[2][10] ), .IN2(n5693), .Q(n5264) );
  AND2X1 U7522 ( .IN1(\decodedPacket[2][11] ), .IN2(n5693), .Q(n5265) );
  INVX0 U7523 ( .INP(\decodedPacket[2][97] ), .ZN(n6114) );
  INVX0 U7524 ( .INP(\decodedPacket[2][79] ), .ZN(n6103) );
  INVX0 U7525 ( .INP(\decodedPacket[2][80] ), .ZN(n6104) );
  INVX0 U7526 ( .INP(\decodedPacket[2][81] ), .ZN(n6105) );
  INVX0 U7527 ( .INP(\decodedPacket[2][82] ), .ZN(n6106) );
  INVX0 U7528 ( .INP(\decodedPacket[2][72] ), .ZN(n6085) );
  INVX0 U7529 ( .INP(\decodedPacket[2][70] ), .ZN(n6043) );
  INVX0 U7530 ( .INP(\decodedPacket[2][115] ), .ZN(n6039) );
  INVX0 U7531 ( .INP(\decodedPacket[2][103] ), .ZN(n6003) );
  INVX0 U7532 ( .INP(\decodedPacket[2][69] ), .ZN(n6084) );
  INVX0 U7533 ( .INP(\decodedPacket[2][99] ), .ZN(n5999) );
  INVX0 U7534 ( .INP(\decodedPacket[2][100] ), .ZN(n6006) );
  INVX0 U7535 ( .INP(\decodedPacket[2][101] ), .ZN(n6005) );
  INVX0 U7536 ( .INP(\decodedPacket[2][102] ), .ZN(n6004) );
  INVX0 U7537 ( .INP(\decodedPacket[2][104] ), .ZN(n6002) );
  INVX0 U7538 ( .INP(\decodedPacket[2][105] ), .ZN(n6001) );
  INVX0 U7539 ( .INP(\decodedPacket[2][106] ), .ZN(n6000) );
  INVX0 U7540 ( .INP(fs2Ready_i), .ZN(n5266) );
  NAND2X1 U7541 ( .IN1(\decodedPacket[0][5] ), .IN2(n5588), .QN(n2488) );
  NAND2X1 U7542 ( .IN1(\decodedPacket[0][6] ), .IN2(n5588), .QN(n2482) );
  NAND2X1 U7543 ( .IN1(\decodedPacket[0][7] ), .IN2(n5588), .QN(n2476) );
  NAND2X1 U7544 ( .IN1(\decodedPacket[0][8] ), .IN2(n5588), .QN(n2470) );
  NAND2X1 U7545 ( .IN1(\decodedPacket[0][9] ), .IN2(n5588), .QN(n2464) );
  NAND2X1 U7546 ( .IN1(\decodedPacket[0][10] ), .IN2(n5588), .QN(n2458) );
  NAND2X1 U7547 ( .IN1(\decodedPacket[0][11] ), .IN2(n5588), .QN(n2452) );
  NAND2X1 U7548 ( .IN1(\decodedPacket[0][12] ), .IN2(n5588), .QN(n2446) );
  NAND2X1 U7549 ( .IN1(\decodedPacket[0][13] ), .IN2(n5588), .QN(n2440) );
  NAND2X1 U7550 ( .IN1(\decodedPacket[0][14] ), .IN2(n5588), .QN(n2434) );
  NAND2X1 U7551 ( .IN1(\decodedPacket[0][15] ), .IN2(n5587), .QN(n2428) );
  NAND2X1 U7552 ( .IN1(\decodedPacket[0][16] ), .IN2(n5587), .QN(n2422) );
  NAND2X1 U7553 ( .IN1(\decodedPacket[0][17] ), .IN2(n5587), .QN(n2416) );
  NAND2X1 U7554 ( .IN1(\decodedPacket[0][18] ), .IN2(n5587), .QN(n2410) );
  NAND2X1 U7555 ( .IN1(\decodedPacket[0][19] ), .IN2(n5587), .QN(n2404) );
  NAND2X1 U7556 ( .IN1(\decodedPacket[0][20] ), .IN2(n5587), .QN(n2398) );
  NAND2X1 U7557 ( .IN1(\decodedPacket[0][21] ), .IN2(n5587), .QN(n2392) );
  NAND2X1 U7558 ( .IN1(\decodedPacket[0][22] ), .IN2(n5587), .QN(n2386) );
  NAND2X1 U7559 ( .IN1(\decodedPacket[0][23] ), .IN2(n5587), .QN(n2380) );
  NAND2X1 U7560 ( .IN1(\decodedPacket[0][24] ), .IN2(n5587), .QN(n2374) );
  NAND2X1 U7561 ( .IN1(\decodedPacket[0][25] ), .IN2(n5587), .QN(n2368) );
  NAND2X1 U7562 ( .IN1(\decodedPacket[0][26] ), .IN2(n5587), .QN(n2362) );
  NAND2X1 U7563 ( .IN1(\decodedPacket[0][27] ), .IN2(n5586), .QN(n2356) );
  NAND2X1 U7564 ( .IN1(\decodedPacket[0][28] ), .IN2(n5586), .QN(n2350) );
  NAND2X1 U7565 ( .IN1(\decodedPacket[0][29] ), .IN2(n5586), .QN(n2344) );
  NAND2X1 U7566 ( .IN1(\decodedPacket[0][30] ), .IN2(n5586), .QN(n2338) );
  NAND2X1 U7567 ( .IN1(\decodedPacket[0][31] ), .IN2(n5586), .QN(n2332) );
  NAND2X1 U7568 ( .IN1(\decodedPacket[0][32] ), .IN2(n5586), .QN(n2326) );
  NAND2X1 U7569 ( .IN1(\decodedPacket[0][33] ), .IN2(n5586), .QN(n2320) );
  NAND2X1 U7570 ( .IN1(\decodedPacket[0][34] ), .IN2(n5586), .QN(n2314) );
  NAND2X1 U7571 ( .IN1(\decodedPacket[0][35] ), .IN2(n5586), .QN(n2308) );
  NAND2X1 U7572 ( .IN1(\decodedPacket[0][36] ), .IN2(n5586), .QN(n2302) );
  INVX0 U7573 ( .INP(\decodedPacket[4][12] ), .ZN(n6190) );
  INVX0 U7574 ( .INP(\decodedPacket[4][13] ), .ZN(n6189) );
  INVX0 U7575 ( .INP(\decodedPacket[4][14] ), .ZN(n6188) );
  INVX0 U7576 ( .INP(\decodedPacket[4][15] ), .ZN(n6187) );
  INVX0 U7577 ( .INP(\decodedPacket[4][16] ), .ZN(n6186) );
  INVX0 U7578 ( .INP(\decodedPacket[4][17] ), .ZN(n6185) );
  INVX0 U7579 ( .INP(\decodedPacket[4][18] ), .ZN(n6184) );
  INVX0 U7580 ( .INP(\decodedPacket[4][19] ), .ZN(n6183) );
  INVX0 U7581 ( .INP(\decodedPacket[4][20] ), .ZN(n6182) );
  INVX0 U7582 ( .INP(\decodedPacket[4][5] ), .ZN(n6165) );
  INVX0 U7583 ( .INP(\decodedPacket[4][6] ), .ZN(n6164) );
  INVX0 U7584 ( .INP(\decodedPacket[4][7] ), .ZN(n6163) );
  INVX0 U7585 ( .INP(\decodedPacket[4][8] ), .ZN(n6162) );
  INVX0 U7586 ( .INP(\decodedPacket[4][9] ), .ZN(n6161) );
  INVX0 U7587 ( .INP(\decodedPacket[4][10] ), .ZN(n6192) );
  INVX0 U7588 ( .INP(\decodedPacket[4][11] ), .ZN(n6191) );
  INVX0 U7589 ( .INP(\decodedPacket[4][21] ), .ZN(n6181) );
  INVX0 U7590 ( .INP(\decodedPacket[4][22] ), .ZN(n6180) );
  INVX0 U7591 ( .INP(\decodedPacket[4][23] ), .ZN(n6179) );
  INVX0 U7592 ( .INP(\decodedPacket[4][24] ), .ZN(n6178) );
  INVX0 U7593 ( .INP(\decodedPacket[4][25] ), .ZN(n6177) );
  INVX0 U7594 ( .INP(\decodedPacket[4][26] ), .ZN(n6176) );
  INVX0 U7595 ( .INP(\decodedPacket[4][27] ), .ZN(n6175) );
  INVX0 U7596 ( .INP(\decodedPacket[4][28] ), .ZN(n6174) );
  INVX0 U7597 ( .INP(\decodedPacket[4][29] ), .ZN(n6173) );
  INVX0 U7598 ( .INP(\decodedPacket[4][30] ), .ZN(n6172) );
  INVX0 U7599 ( .INP(\decodedPacket[4][31] ), .ZN(n6171) );
  INVX0 U7600 ( .INP(\decodedPacket[4][32] ), .ZN(n6170) );
  INVX0 U7601 ( .INP(\decodedPacket[4][33] ), .ZN(n6169) );
  INVX0 U7602 ( .INP(\decodedPacket[4][34] ), .ZN(n6168) );
  INVX0 U7603 ( .INP(\decodedPacket[4][35] ), .ZN(n6167) );
  INVX0 U7604 ( .INP(\decodedPacket[4][36] ), .ZN(n6166) );
  INVX0 U7605 ( .INP(\decodedPacket[4][112] ), .ZN(n6213) );
  INVX0 U7606 ( .INP(\decodedPacket[4][113] ), .ZN(n6214) );
  INVX0 U7607 ( .INP(\decodedPacket[4][114] ), .ZN(n6215) );
  INVX0 U7608 ( .INP(\decodedPacket[6][112] ), .ZN(n6367) );
  INVX0 U7609 ( .INP(\decodedPacket[6][113] ), .ZN(n6368) );
  INVX0 U7610 ( .INP(\decodedPacket[6][114] ), .ZN(n6369) );
  INVX0 U7611 ( .INP(\decodedPacket[4][97] ), .ZN(n6268) );
  INVX0 U7612 ( .INP(\decodedPacket[6][97] ), .ZN(n6422) );
  INVX0 U7613 ( .INP(\decodedPacket[4][79] ), .ZN(n6257) );
  INVX0 U7614 ( .INP(\decodedPacket[4][80] ), .ZN(n6258) );
  INVX0 U7615 ( .INP(\decodedPacket[4][81] ), .ZN(n6259) );
  INVX0 U7616 ( .INP(\decodedPacket[4][82] ), .ZN(n6260) );
  INVX0 U7617 ( .INP(\decodedPacket[6][79] ), .ZN(n6411) );
  INVX0 U7618 ( .INP(\decodedPacket[6][80] ), .ZN(n6412) );
  INVX0 U7619 ( .INP(\decodedPacket[6][81] ), .ZN(n6413) );
  INVX0 U7620 ( .INP(\decodedPacket[6][82] ), .ZN(n6414) );
  INVX0 U7621 ( .INP(\decodedPacket[6][12] ), .ZN(n6344) );
  INVX0 U7622 ( .INP(\decodedPacket[6][13] ), .ZN(n6343) );
  INVX0 U7623 ( .INP(\decodedPacket[6][14] ), .ZN(n6342) );
  INVX0 U7624 ( .INP(\decodedPacket[6][15] ), .ZN(n6341) );
  INVX0 U7625 ( .INP(\decodedPacket[6][16] ), .ZN(n6340) );
  INVX0 U7626 ( .INP(\decodedPacket[6][5] ), .ZN(n6319) );
  INVX0 U7627 ( .INP(\decodedPacket[6][6] ), .ZN(n6318) );
  INVX0 U7628 ( .INP(\decodedPacket[6][7] ), .ZN(n6317) );
  INVX0 U7629 ( .INP(\decodedPacket[6][8] ), .ZN(n6316) );
  INVX0 U7630 ( .INP(\decodedPacket[6][9] ), .ZN(n6315) );
  INVX0 U7631 ( .INP(\decodedPacket[6][10] ), .ZN(n6346) );
  INVX0 U7632 ( .INP(\decodedPacket[6][11] ), .ZN(n6345) );
  INVX0 U7633 ( .INP(\decodedPacket[6][17] ), .ZN(n6339) );
  INVX0 U7634 ( .INP(\decodedPacket[6][18] ), .ZN(n6338) );
  INVX0 U7635 ( .INP(\decodedPacket[6][19] ), .ZN(n6337) );
  INVX0 U7636 ( .INP(\decodedPacket[6][20] ), .ZN(n6336) );
  INVX0 U7637 ( .INP(\decodedPacket[6][21] ), .ZN(n6335) );
  INVX0 U7638 ( .INP(\decodedPacket[6][22] ), .ZN(n6334) );
  INVX0 U7639 ( .INP(\decodedPacket[6][23] ), .ZN(n6333) );
  INVX0 U7640 ( .INP(\decodedPacket[6][24] ), .ZN(n6332) );
  INVX0 U7641 ( .INP(\decodedPacket[6][25] ), .ZN(n6331) );
  INVX0 U7642 ( .INP(\decodedPacket[6][26] ), .ZN(n6330) );
  INVX0 U7643 ( .INP(\decodedPacket[6][27] ), .ZN(n6329) );
  INVX0 U7644 ( .INP(\decodedPacket[6][28] ), .ZN(n6328) );
  INVX0 U7645 ( .INP(\decodedPacket[6][29] ), .ZN(n6327) );
  INVX0 U7646 ( .INP(\decodedPacket[6][30] ), .ZN(n6326) );
  INVX0 U7647 ( .INP(\decodedPacket[4][72] ), .ZN(n6239) );
  INVX0 U7648 ( .INP(\decodedPacket[6][72] ), .ZN(n6393) );
  INVX0 U7649 ( .INP(\decodedPacket[4][70] ), .ZN(n6197) );
  INVX0 U7650 ( .INP(\decodedPacket[6][70] ), .ZN(n6351) );
  INVX0 U7651 ( .INP(\decodedPacket[3][90] ), .ZN(n6077) );
  INVX0 U7652 ( .INP(\decodedPacket[3][86] ), .ZN(n6081) );
  INVX0 U7653 ( .INP(\decodedPacket[3][87] ), .ZN(n6080) );
  INVX0 U7654 ( .INP(\decodedPacket[3][88] ), .ZN(n6079) );
  INVX0 U7655 ( .INP(\decodedPacket[3][89] ), .ZN(n6078) );
  INVX0 U7656 ( .INP(\decodedPacket[3][85] ), .ZN(n6082) );
  INVX0 U7657 ( .INP(\decodedPacket[5][90] ), .ZN(n6231) );
  INVX0 U7658 ( .INP(\decodedPacket[5][86] ), .ZN(n6235) );
  INVX0 U7659 ( .INP(\decodedPacket[5][87] ), .ZN(n6234) );
  INVX0 U7660 ( .INP(\decodedPacket[5][88] ), .ZN(n6233) );
  INVX0 U7661 ( .INP(\decodedPacket[5][89] ), .ZN(n6232) );
  INVX0 U7662 ( .INP(\decodedPacket[5][85] ), .ZN(n6236) );
  INVX0 U7663 ( .INP(\decodedPacket[4][115] ), .ZN(n6193) );
  INVX0 U7664 ( .INP(\decodedPacket[6][115] ), .ZN(n6347) );
  INVX0 U7665 ( .INP(\decodedPacket[4][103] ), .ZN(n6157) );
  INVX0 U7666 ( .INP(\decodedPacket[6][103] ), .ZN(n6311) );
  INVX0 U7667 ( .INP(\decodedPacket[4][69] ), .ZN(n6238) );
  INVX0 U7668 ( .INP(\decodedPacket[6][69] ), .ZN(n6392) );
  INVX0 U7669 ( .INP(\decodedPacket[4][99] ), .ZN(n6153) );
  INVX0 U7670 ( .INP(\decodedPacket[4][100] ), .ZN(n6160) );
  INVX0 U7671 ( .INP(\decodedPacket[4][101] ), .ZN(n6159) );
  INVX0 U7672 ( .INP(\decodedPacket[4][102] ), .ZN(n6158) );
  INVX0 U7673 ( .INP(\decodedPacket[4][104] ), .ZN(n6156) );
  INVX0 U7674 ( .INP(\decodedPacket[4][105] ), .ZN(n6155) );
  INVX0 U7675 ( .INP(\decodedPacket[4][106] ), .ZN(n6154) );
  INVX0 U7676 ( .INP(\decodedPacket[6][99] ), .ZN(n6307) );
  INVX0 U7677 ( .INP(\decodedPacket[6][100] ), .ZN(n6314) );
  INVX0 U7678 ( .INP(\decodedPacket[6][101] ), .ZN(n6313) );
  INVX0 U7679 ( .INP(\decodedPacket[6][102] ), .ZN(n6312) );
  INVX0 U7680 ( .INP(\decodedPacket[6][104] ), .ZN(n6310) );
  INVX0 U7681 ( .INP(\decodedPacket[6][105] ), .ZN(n6309) );
  INVX0 U7682 ( .INP(\decodedPacket[6][106] ), .ZN(n6308) );
  INVX0 U7683 ( .INP(\decodedPacket[6][31] ), .ZN(n6325) );
  INVX0 U7684 ( .INP(\decodedPacket[6][32] ), .ZN(n6324) );
  INVX0 U7685 ( .INP(\decodedPacket[6][33] ), .ZN(n6323) );
  INVX0 U7686 ( .INP(\decodedPacket[6][34] ), .ZN(n6322) );
  INVX0 U7687 ( .INP(\decodedPacket[6][35] ), .ZN(n6321) );
  INVX0 U7688 ( .INP(\decodedPacket[6][36] ), .ZN(n6320) );
  INVX0 U7689 ( .INP(\decodedPacket[6][0] ), .ZN(n6459) );
  INVX0 U7690 ( .INP(\decodedPacket[6][1] ), .ZN(n6458) );
  INVX0 U7691 ( .INP(\decodedPacket[6][38] ), .ZN(n6453) );
  INVX0 U7692 ( .INP(\decodedPacket[6][39] ), .ZN(n6452) );
  INVX0 U7693 ( .INP(\decodedPacket[6][40] ), .ZN(n6451) );
  INVX0 U7694 ( .INP(\decodedPacket[6][41] ), .ZN(n6450) );
  INVX0 U7695 ( .INP(\decodedPacket[6][42] ), .ZN(n6449) );
  INVX0 U7696 ( .INP(\decodedPacket[6][43] ), .ZN(n6448) );
  INVX0 U7697 ( .INP(\decodedPacket[6][44] ), .ZN(n6447) );
  INVX0 U7698 ( .INP(\decodedPacket[3][99] ), .ZN(n6067) );
  INVX0 U7699 ( .INP(\decodedPacket[3][100] ), .ZN(n5951) );
  INVX0 U7700 ( .INP(\decodedPacket[3][101] ), .ZN(n5950) );
  INVX0 U7701 ( .INP(\decodedPacket[3][102] ), .ZN(n5949) );
  INVX0 U7702 ( .INP(\decodedPacket[3][103] ), .ZN(n5948) );
  INVX0 U7703 ( .INP(\decodedPacket[3][104] ), .ZN(n5947) );
  INVX0 U7704 ( .INP(\decodedPacket[3][105] ), .ZN(n5946) );
  INVX0 U7705 ( .INP(\decodedPacket[3][106] ), .ZN(n5945) );
  INVX0 U7706 ( .INP(\decodedPacket[3][107] ), .ZN(n5944) );
  INVX0 U7707 ( .INP(\decodedPacket[3][108] ), .ZN(n5943) );
  INVX0 U7708 ( .INP(\decodedPacket[3][109] ), .ZN(n5942) );
  INVX0 U7709 ( .INP(\decodedPacket[3][110] ), .ZN(n5941) );
  INVX0 U7710 ( .INP(\decodedPacket[3][111] ), .ZN(n5940) );
  INVX0 U7711 ( .INP(\decodedPacket[3][112] ), .ZN(n5939) );
  INVX0 U7712 ( .INP(\decodedPacket[3][113] ), .ZN(n5938) );
  INVX0 U7713 ( .INP(\decodedPacket[3][79] ), .ZN(n6101) );
  INVX0 U7714 ( .INP(\decodedPacket[3][80] ), .ZN(n6100) );
  INVX0 U7715 ( .INP(\decodedPacket[3][81] ), .ZN(n6099) );
  INVX0 U7716 ( .INP(\decodedPacket[3][82] ), .ZN(n6098) );
  INVX0 U7717 ( .INP(\decodedPacket[5][99] ), .ZN(n6221) );
  INVX0 U7718 ( .INP(\decodedPacket[5][100] ), .ZN(n5966) );
  INVX0 U7719 ( .INP(\decodedPacket[5][101] ), .ZN(n5965) );
  INVX0 U7720 ( .INP(\decodedPacket[5][102] ), .ZN(n5964) );
  INVX0 U7721 ( .INP(\decodedPacket[5][103] ), .ZN(n5963) );
  INVX0 U7722 ( .INP(\decodedPacket[5][104] ), .ZN(n5962) );
  INVX0 U7723 ( .INP(\decodedPacket[5][105] ), .ZN(n5961) );
  INVX0 U7724 ( .INP(\decodedPacket[5][106] ), .ZN(n5960) );
  INVX0 U7725 ( .INP(\decodedPacket[5][107] ), .ZN(n5959) );
  INVX0 U7726 ( .INP(\decodedPacket[5][108] ), .ZN(n5958) );
  INVX0 U7727 ( .INP(\decodedPacket[5][109] ), .ZN(n5957) );
  INVX0 U7728 ( .INP(\decodedPacket[5][110] ), .ZN(n5956) );
  INVX0 U7729 ( .INP(\decodedPacket[5][111] ), .ZN(n5955) );
  INVX0 U7730 ( .INP(\decodedPacket[5][112] ), .ZN(n5954) );
  INVX0 U7731 ( .INP(\decodedPacket[5][113] ), .ZN(n5953) );
  INVX0 U7732 ( .INP(\decodedPacket[5][79] ), .ZN(n6255) );
  INVX0 U7733 ( .INP(\decodedPacket[5][80] ), .ZN(n6254) );
  INVX0 U7734 ( .INP(\decodedPacket[5][81] ), .ZN(n6253) );
  INVX0 U7735 ( .INP(\decodedPacket[5][82] ), .ZN(n6252) );
  INVX0 U7736 ( .INP(\decodedPacket[4][0] ), .ZN(n6305) );
  INVX0 U7737 ( .INP(\decodedPacket[4][1] ), .ZN(n6304) );
  INVX0 U7738 ( .INP(\decodedPacket[4][2] ), .ZN(n6303) );
  INVX0 U7739 ( .INP(\decodedPacket[4][3] ), .ZN(n6302) );
  INVX0 U7740 ( .INP(\decodedPacket[4][4] ), .ZN(n6301) );
  INVX0 U7741 ( .INP(\decodedPacket[4][37] ), .ZN(n6300) );
  INVX0 U7742 ( .INP(\decodedPacket[4][38] ), .ZN(n6299) );
  INVX0 U7743 ( .INP(\decodedPacket[4][39] ), .ZN(n6298) );
  INVX0 U7744 ( .INP(\decodedPacket[4][40] ), .ZN(n6297) );
  INVX0 U7745 ( .INP(\decodedPacket[4][41] ), .ZN(n6296) );
  INVX0 U7746 ( .INP(\decodedPacket[4][42] ), .ZN(n6295) );
  INVX0 U7747 ( .INP(\decodedPacket[4][43] ), .ZN(n6294) );
  INVX0 U7748 ( .INP(\decodedPacket[4][44] ), .ZN(n6293) );
  INVX0 U7749 ( .INP(\decodedPacket[4][45] ), .ZN(n6292) );
  INVX0 U7750 ( .INP(\decodedPacket[4][46] ), .ZN(n6291) );
  INVX0 U7751 ( .INP(\decodedPacket[4][47] ), .ZN(n6290) );
  INVX0 U7752 ( .INP(\decodedPacket[4][48] ), .ZN(n6289) );
  INVX0 U7753 ( .INP(\decodedPacket[4][49] ), .ZN(n6288) );
  INVX0 U7754 ( .INP(\decodedPacket[4][50] ), .ZN(n6287) );
  INVX0 U7755 ( .INP(\decodedPacket[4][51] ), .ZN(n6286) );
  INVX0 U7756 ( .INP(\decodedPacket[4][52] ), .ZN(n6285) );
  INVX0 U7757 ( .INP(\decodedPacket[4][53] ), .ZN(n6284) );
  INVX0 U7758 ( .INP(\decodedPacket[4][54] ), .ZN(n6283) );
  INVX0 U7759 ( .INP(\decodedPacket[4][55] ), .ZN(n6282) );
  INVX0 U7760 ( .INP(\decodedPacket[4][56] ), .ZN(n6281) );
  INVX0 U7761 ( .INP(\decodedPacket[4][57] ), .ZN(n6280) );
  INVX0 U7762 ( .INP(\decodedPacket[4][58] ), .ZN(n6279) );
  INVX0 U7763 ( .INP(\decodedPacket[4][59] ), .ZN(n6278) );
  INVX0 U7764 ( .INP(\decodedPacket[4][60] ), .ZN(n6277) );
  INVX0 U7765 ( .INP(\decodedPacket[4][61] ), .ZN(n6276) );
  INVX0 U7766 ( .INP(\decodedPacket[4][62] ), .ZN(n6275) );
  INVX0 U7767 ( .INP(\decodedPacket[4][63] ), .ZN(n6274) );
  INVX0 U7768 ( .INP(\decodedPacket[4][64] ), .ZN(n6273) );
  INVX0 U7769 ( .INP(\decodedPacket[4][65] ), .ZN(n6272) );
  INVX0 U7770 ( .INP(\decodedPacket[4][66] ), .ZN(n6271) );
  INVX0 U7771 ( .INP(\decodedPacket[4][67] ), .ZN(n6270) );
  INVX0 U7772 ( .INP(\decodedPacket[4][68] ), .ZN(n6269) );
  INVX0 U7773 ( .INP(\decodedPacket[6][45] ), .ZN(n6446) );
  INVX0 U7774 ( .INP(\decodedPacket[6][46] ), .ZN(n6445) );
  INVX0 U7775 ( .INP(\decodedPacket[6][47] ), .ZN(n6444) );
  INVX0 U7776 ( .INP(\decodedPacket[6][48] ), .ZN(n6443) );
  INVX0 U7777 ( .INP(\decodedPacket[6][49] ), .ZN(n6442) );
  INVX0 U7778 ( .INP(\decodedPacket[6][50] ), .ZN(n6441) );
  INVX0 U7779 ( .INP(\decodedPacket[6][51] ), .ZN(n6440) );
  INVX0 U7780 ( .INP(\decodedPacket[6][52] ), .ZN(n6439) );
  INVX0 U7781 ( .INP(\decodedPacket[6][53] ), .ZN(n6438) );
  INVX0 U7782 ( .INP(\decodedPacket[6][54] ), .ZN(n6437) );
  INVX0 U7783 ( .INP(\decodedPacket[6][55] ), .ZN(n6436) );
  INVX0 U7784 ( .INP(\decodedPacket[6][56] ), .ZN(n6435) );
  INVX0 U7785 ( .INP(\decodedPacket[6][57] ), .ZN(n6434) );
  INVX0 U7786 ( .INP(\decodedPacket[6][58] ), .ZN(n6433) );
  INVX0 U7787 ( .INP(\decodedPacket[6][59] ), .ZN(n6432) );
  INVX0 U7788 ( .INP(\decodedPacket[6][60] ), .ZN(n6431) );
  INVX0 U7789 ( .INP(\decodedPacket[6][61] ), .ZN(n6430) );
  INVX0 U7790 ( .INP(\decodedPacket[6][62] ), .ZN(n6429) );
  INVX0 U7791 ( .INP(\decodedPacket[6][63] ), .ZN(n6428) );
  INVX0 U7792 ( .INP(\decodedPacket[6][64] ), .ZN(n6427) );
  INVX0 U7793 ( .INP(\decodedPacket[6][65] ), .ZN(n6426) );
  INVX0 U7794 ( .INP(\decodedPacket[6][66] ), .ZN(n6425) );
  INVX0 U7795 ( .INP(\decodedPacket[6][67] ), .ZN(n6424) );
  INVX0 U7796 ( .INP(\decodedPacket[6][68] ), .ZN(n6423) );
  INVX0 U7797 ( .INP(\decodedPacket[3][0] ), .ZN(n6151) );
  INVX0 U7798 ( .INP(\decodedPacket[3][1] ), .ZN(n6150) );
  INVX0 U7799 ( .INP(\decodedPacket[3][2] ), .ZN(n6149) );
  INVX0 U7800 ( .INP(\decodedPacket[3][3] ), .ZN(n6148) );
  INVX0 U7801 ( .INP(\decodedPacket[3][4] ), .ZN(n6147) );
  INVX0 U7802 ( .INP(\decodedPacket[3][37] ), .ZN(n6146) );
  INVX0 U7803 ( .INP(\decodedPacket[3][38] ), .ZN(n6145) );
  INVX0 U7804 ( .INP(\decodedPacket[3][39] ), .ZN(n6144) );
  INVX0 U7805 ( .INP(\decodedPacket[3][40] ), .ZN(n6143) );
  INVX0 U7806 ( .INP(\decodedPacket[3][41] ), .ZN(n6142) );
  INVX0 U7807 ( .INP(\decodedPacket[3][42] ), .ZN(n6141) );
  INVX0 U7808 ( .INP(\decodedPacket[3][43] ), .ZN(n6140) );
  INVX0 U7809 ( .INP(\decodedPacket[3][44] ), .ZN(n6139) );
  INVX0 U7810 ( .INP(\decodedPacket[3][45] ), .ZN(n6138) );
  INVX0 U7811 ( .INP(\decodedPacket[3][46] ), .ZN(n6137) );
  INVX0 U7812 ( .INP(\decodedPacket[3][47] ), .ZN(n6136) );
  INVX0 U7813 ( .INP(\decodedPacket[3][48] ), .ZN(n6135) );
  INVX0 U7814 ( .INP(\decodedPacket[3][49] ), .ZN(n6134) );
  INVX0 U7815 ( .INP(\decodedPacket[3][50] ), .ZN(n6133) );
  INVX0 U7816 ( .INP(\decodedPacket[3][51] ), .ZN(n6132) );
  INVX0 U7817 ( .INP(\decodedPacket[3][52] ), .ZN(n6131) );
  INVX0 U7818 ( .INP(\decodedPacket[3][53] ), .ZN(n6130) );
  INVX0 U7819 ( .INP(\decodedPacket[3][54] ), .ZN(n6129) );
  INVX0 U7820 ( .INP(\decodedPacket[3][55] ), .ZN(n6128) );
  INVX0 U7821 ( .INP(\decodedPacket[3][56] ), .ZN(n6127) );
  INVX0 U7822 ( .INP(\decodedPacket[3][57] ), .ZN(n6126) );
  INVX0 U7823 ( .INP(\decodedPacket[3][58] ), .ZN(n6125) );
  INVX0 U7824 ( .INP(\decodedPacket[3][59] ), .ZN(n6124) );
  INVX0 U7825 ( .INP(\decodedPacket[3][60] ), .ZN(n6123) );
  INVX0 U7826 ( .INP(\decodedPacket[3][61] ), .ZN(n6122) );
  INVX0 U7827 ( .INP(\decodedPacket[3][62] ), .ZN(n6121) );
  INVX0 U7828 ( .INP(\decodedPacket[3][63] ), .ZN(n6120) );
  INVX0 U7829 ( .INP(\decodedPacket[3][64] ), .ZN(n6119) );
  INVX0 U7830 ( .INP(\decodedPacket[3][65] ), .ZN(n6118) );
  INVX0 U7831 ( .INP(\decodedPacket[3][66] ), .ZN(n6117) );
  INVX0 U7832 ( .INP(\decodedPacket[3][67] ), .ZN(n6116) );
  INVX0 U7833 ( .INP(\decodedPacket[3][68] ), .ZN(n6115) );
  INVX0 U7834 ( .INP(\decodedPacket[7][90] ), .ZN(n6385) );
  INVX0 U7835 ( .INP(\decodedPacket[7][86] ), .ZN(n6389) );
  INVX0 U7836 ( .INP(\decodedPacket[7][87] ), .ZN(n6388) );
  INVX0 U7837 ( .INP(\decodedPacket[7][88] ), .ZN(n6387) );
  INVX0 U7838 ( .INP(\decodedPacket[7][89] ), .ZN(n6386) );
  INVX0 U7839 ( .INP(\decodedPacket[7][85] ), .ZN(n6390) );
  INVX0 U7840 ( .INP(\decodedPacket[7][2] ), .ZN(n6457) );
  INVX0 U7841 ( .INP(\decodedPacket[7][3] ), .ZN(n6456) );
  INVX0 U7842 ( .INP(\decodedPacket[7][4] ), .ZN(n6455) );
  INVX0 U7843 ( .INP(\decodedPacket[7][37] ), .ZN(n6454) );
  INVX0 U7844 ( .INP(\decodedPacket[7][99] ), .ZN(n6375) );
  INVX0 U7845 ( .INP(\decodedPacket[7][100] ), .ZN(n5981) );
  INVX0 U7846 ( .INP(\decodedPacket[7][101] ), .ZN(n5980) );
  INVX0 U7847 ( .INP(\decodedPacket[7][102] ), .ZN(n5979) );
  INVX0 U7848 ( .INP(\decodedPacket[7][103] ), .ZN(n5978) );
  INVX0 U7849 ( .INP(\decodedPacket[7][104] ), .ZN(n5977) );
  INVX0 U7850 ( .INP(\decodedPacket[7][105] ), .ZN(n5976) );
  INVX0 U7851 ( .INP(\decodedPacket[7][106] ), .ZN(n5975) );
  INVX0 U7852 ( .INP(\decodedPacket[7][107] ), .ZN(n5974) );
  INVX0 U7853 ( .INP(\decodedPacket[7][108] ), .ZN(n5973) );
  INVX0 U7854 ( .INP(\decodedPacket[7][109] ), .ZN(n5972) );
  INVX0 U7855 ( .INP(\decodedPacket[7][110] ), .ZN(n5971) );
  INVX0 U7856 ( .INP(\decodedPacket[7][111] ), .ZN(n5970) );
  INVX0 U7857 ( .INP(\decodedPacket[7][112] ), .ZN(n5969) );
  INVX0 U7858 ( .INP(\decodedPacket[7][113] ), .ZN(n5968) );
  INVX0 U7859 ( .INP(\decodedPacket[7][79] ), .ZN(n6409) );
  INVX0 U7860 ( .INP(\decodedPacket[7][80] ), .ZN(n6408) );
  INVX0 U7861 ( .INP(\decodedPacket[7][81] ), .ZN(n6407) );
  INVX0 U7862 ( .INP(\decodedPacket[7][82] ), .ZN(n6406) );
  INVX0 U7863 ( .INP(n5266), .ZN(decodeReady_o) );
  INVX0 U7896 ( .INP(n5282), .ZN(n5276) );
  INVX0 U7897 ( .INP(n5282), .ZN(n5277) );
  INVX0 U7898 ( .INP(n5282), .ZN(n5278) );
  INVX0 U7899 ( .INP(n5282), .ZN(n5279) );
  INVX0 U7900 ( .INP(n5282), .ZN(n5280) );
  INVX0 U7901 ( .INP(n5282), .ZN(n5281) );
  NBUFFX2 U7902 ( .INP(n4076), .Z(n5284) );
  NBUFFX2 U7903 ( .INP(n4076), .Z(n5285) );
  INVX0 U7904 ( .INP(n5296), .ZN(n5286) );
  INVX0 U7905 ( .INP(n5296), .ZN(n5287) );
  INVX0 U7906 ( .INP(n5296), .ZN(n5288) );
  INVX0 U7907 ( .INP(n5296), .ZN(n5289) );
  INVX0 U7908 ( .INP(n5296), .ZN(n5290) );
  INVX0 U7909 ( .INP(n5296), .ZN(n5291) );
  INVX0 U7910 ( .INP(n5296), .ZN(n5292) );
  INVX0 U7911 ( .INP(n5296), .ZN(n5293) );
  INVX0 U7912 ( .INP(n5296), .ZN(n5294) );
  INVX0 U7913 ( .INP(n5296), .ZN(n5295) );
  NBUFFX2 U7914 ( .INP(n4076), .Z(n5296) );
  NBUFFX2 U7915 ( .INP(n5284), .Z(n5297) );
  NBUFFX2 U7916 ( .INP(n5285), .Z(n5298) );
  NBUFFX2 U7917 ( .INP(n5284), .Z(n5299) );
  NBUFFX2 U7918 ( .INP(n5284), .Z(n5300) );
  NBUFFX2 U7919 ( .INP(n5285), .Z(n5301) );
  NBUFFX2 U7920 ( .INP(n5285), .Z(n5302) );
  NBUFFX2 U7921 ( .INP(n5285), .Z(n5303) );
  INVX0 U7922 ( .INP(n5312), .ZN(n5304) );
  INVX0 U7923 ( .INP(n5316), .ZN(n5305) );
  INVX0 U7924 ( .INP(n4916), .ZN(n5306) );
  INVX0 U7925 ( .INP(n5310), .ZN(n5307) );
  INVX0 U7926 ( .INP(n5316), .ZN(n5308) );
  INVX0 U7927 ( .INP(n5313), .ZN(n5309) );
  NBUFFX2 U7928 ( .INP(n4072), .Z(n5318) );
  NBUFFX2 U7929 ( .INP(n4072), .Z(n5319) );
  NBUFFX2 U7930 ( .INP(n4072), .Z(n5320) );
  INVX0 U7931 ( .INP(n5318), .ZN(n5321) );
  INVX0 U7932 ( .INP(n5318), .ZN(n5322) );
  INVX0 U7933 ( .INP(n5318), .ZN(n5323) );
  INVX0 U7934 ( .INP(n5318), .ZN(n5324) );
  INVX0 U7935 ( .INP(n5318), .ZN(n5325) );
  INVX0 U7936 ( .INP(n5318), .ZN(n5326) );
  INVX0 U7937 ( .INP(n5318), .ZN(n5327) );
  INVX0 U7938 ( .INP(n5318), .ZN(n5328) );
  INVX0 U7939 ( .INP(n5320), .ZN(n5329) );
  INVX0 U7940 ( .INP(n5318), .ZN(n5330) );
  NBUFFX2 U7941 ( .INP(n5318), .Z(n5331) );
  NBUFFX2 U7942 ( .INP(n5318), .Z(n5332) );
  NBUFFX2 U7943 ( .INP(n5319), .Z(n5333) );
  NBUFFX2 U7944 ( .INP(n5319), .Z(n5334) );
  NBUFFX2 U7945 ( .INP(n5319), .Z(n5335) );
  NBUFFX2 U7946 ( .INP(n5320), .Z(n5336) );
  NBUFFX2 U7947 ( .INP(n5320), .Z(n5337) );
  INVX0 U7948 ( .INP(n5347), .ZN(n5338) );
  INVX0 U7949 ( .INP(n5344), .ZN(n5339) );
  INVX0 U7950 ( .INP(n4070), .ZN(n5340) );
  INVX0 U7951 ( .INP(n5345), .ZN(n5341) );
  INVX0 U7952 ( .INP(n5346), .ZN(n5342) );
  INVX0 U7953 ( .INP(n3686), .ZN(n5351) );
  INVX0 U7954 ( .INP(n5360), .ZN(n5352) );
  INVX0 U7955 ( .INP(n5359), .ZN(n5353) );
  INVX0 U7956 ( .INP(n5360), .ZN(n5354) );
  INVX0 U7957 ( .INP(n5376), .ZN(n5363) );
  INVX0 U7958 ( .INP(n5376), .ZN(n5364) );
  INVX0 U7959 ( .INP(n5376), .ZN(n5365) );
  INVX0 U7960 ( .INP(n5376), .ZN(n5366) );
  INVX0 U7961 ( .INP(n5376), .ZN(n5367) );
  INVX0 U7962 ( .INP(n5376), .ZN(n5368) );
  NBUFFX2 U7963 ( .INP(n5374), .Z(n5369) );
  NBUFFX2 U7964 ( .INP(n5375), .Z(n5370) );
  NBUFFX2 U7965 ( .INP(n5374), .Z(n5371) );
  NBUFFX2 U7966 ( .INP(n5375), .Z(n5372) );
  NBUFFX2 U7967 ( .INP(n5374), .Z(n5373) );
  NBUFFX2 U7968 ( .INP(n4911), .Z(n5374) );
  NBUFFX2 U7969 ( .INP(n4911), .Z(n5375) );
  NBUFFX2 U7970 ( .INP(n4911), .Z(n5376) );
  INVX0 U7971 ( .INP(n5396), .ZN(n5377) );
  INVX0 U7972 ( .INP(n5386), .ZN(n5378) );
  INVX0 U7973 ( .INP(n5391), .ZN(n5379) );
  INVX0 U7974 ( .INP(n5390), .ZN(n5380) );
  INVX0 U7975 ( .INP(n5393), .ZN(n5381) );
  INVX0 U7976 ( .INP(n5388), .ZN(n5382) );
  INVX0 U7977 ( .INP(n5391), .ZN(n5383) );
  INVX0 U7978 ( .INP(n5388), .ZN(n5384) );
  INVX0 U7979 ( .INP(n5387), .ZN(n5385) );
  INVX0 U7980 ( .INP(n3682), .ZN(n5394) );
  INVX0 U7981 ( .INP(n3682), .ZN(n5395) );
  INVX0 U7982 ( .INP(n3682), .ZN(n5396) );
  INVX0 U7983 ( .INP(n5407), .ZN(n5399) );
  INVX0 U7984 ( .INP(n5398), .ZN(n5400) );
  INVX0 U7985 ( .INP(n3680), .ZN(n5401) );
  INVX0 U7986 ( .INP(n5397), .ZN(n5402) );
  INVX0 U7987 ( .INP(n5409), .ZN(n5403) );
  INVX0 U7988 ( .INP(n3302), .ZN(n5410) );
  INVX0 U7989 ( .INP(n5417), .ZN(n5411) );
  INVX0 U7990 ( .INP(n5417), .ZN(n5412) );
  INVX0 U7991 ( .INP(n5415), .ZN(n5413) );
  INVX0 U7992 ( .INP(n5435), .ZN(n5422) );
  INVX0 U7993 ( .INP(n5435), .ZN(n5423) );
  INVX0 U7994 ( .INP(n5435), .ZN(n5424) );
  INVX0 U7995 ( .INP(n5435), .ZN(n5425) );
  INVX0 U7996 ( .INP(n5435), .ZN(n5426) );
  INVX0 U7997 ( .INP(n5435), .ZN(n5427) );
  NBUFFX2 U7998 ( .INP(n5433), .Z(n5428) );
  NBUFFX2 U7999 ( .INP(n5434), .Z(n5429) );
  NBUFFX2 U8000 ( .INP(n5433), .Z(n5430) );
  NBUFFX2 U8001 ( .INP(n5434), .Z(n5431) );
  NBUFFX2 U8002 ( .INP(n5433), .Z(n5432) );
  NBUFFX2 U8003 ( .INP(n4912), .Z(n5433) );
  NBUFFX2 U8004 ( .INP(n4912), .Z(n5434) );
  NBUFFX2 U8005 ( .INP(n4912), .Z(n5435) );
  INVX0 U8006 ( .INP(n5455), .ZN(n5436) );
  INVX0 U8007 ( .INP(n5445), .ZN(n5437) );
  INVX0 U8008 ( .INP(n5450), .ZN(n5438) );
  INVX0 U8009 ( .INP(n5449), .ZN(n5439) );
  INVX0 U8010 ( .INP(n5452), .ZN(n5440) );
  INVX0 U8011 ( .INP(n5447), .ZN(n5441) );
  INVX0 U8012 ( .INP(n5450), .ZN(n5442) );
  INVX0 U8013 ( .INP(n5447), .ZN(n5443) );
  INVX0 U8014 ( .INP(n5446), .ZN(n5444) );
  INVX0 U8015 ( .INP(n3298), .ZN(n5453) );
  INVX0 U8016 ( .INP(n3298), .ZN(n5454) );
  INVX0 U8017 ( .INP(n3298), .ZN(n5455) );
  INVX0 U8018 ( .INP(n5463), .ZN(n5458) );
  INVX0 U8019 ( .INP(n5464), .ZN(n5459) );
  INVX0 U8020 ( .INP(n3296), .ZN(n5460) );
  INVX0 U8021 ( .INP(n5465), .ZN(n5461) );
  INVX0 U8022 ( .INP(n5467), .ZN(n5462) );
  INVX0 U8023 ( .INP(n2918), .ZN(n5469) );
  INVX0 U8024 ( .INP(n5478), .ZN(n5470) );
  INVX0 U8025 ( .INP(n5475), .ZN(n5471) );
  INVX0 U8026 ( .INP(n5478), .ZN(n5472) );
  INVX0 U8027 ( .INP(n5494), .ZN(n5481) );
  INVX0 U8028 ( .INP(n5494), .ZN(n5482) );
  INVX0 U8029 ( .INP(n5494), .ZN(n5483) );
  INVX0 U8030 ( .INP(n5494), .ZN(n5484) );
  INVX0 U8031 ( .INP(n5494), .ZN(n5485) );
  INVX0 U8032 ( .INP(n5494), .ZN(n5486) );
  NBUFFX2 U8033 ( .INP(n5492), .Z(n5487) );
  NBUFFX2 U8034 ( .INP(n5493), .Z(n5488) );
  NBUFFX2 U8035 ( .INP(n5492), .Z(n5489) );
  NBUFFX2 U8036 ( .INP(n5493), .Z(n5490) );
  NBUFFX2 U8037 ( .INP(n5492), .Z(n5491) );
  NBUFFX2 U8038 ( .INP(n4913), .Z(n5492) );
  NBUFFX2 U8039 ( .INP(n4913), .Z(n5493) );
  NBUFFX2 U8040 ( .INP(n4913), .Z(n5494) );
  INVX0 U8041 ( .INP(n5514), .ZN(n5495) );
  INVX0 U8042 ( .INP(n5504), .ZN(n5496) );
  INVX0 U8043 ( .INP(n5509), .ZN(n5497) );
  INVX0 U8044 ( .INP(n5508), .ZN(n5498) );
  INVX0 U8045 ( .INP(n5511), .ZN(n5499) );
  INVX0 U8046 ( .INP(n5506), .ZN(n5500) );
  INVX0 U8047 ( .INP(n5509), .ZN(n5501) );
  INVX0 U8048 ( .INP(n5506), .ZN(n5502) );
  INVX0 U8049 ( .INP(n5505), .ZN(n5503) );
  INVX0 U8050 ( .INP(n2914), .ZN(n5512) );
  INVX0 U8051 ( .INP(n2914), .ZN(n5513) );
  INVX0 U8052 ( .INP(n2914), .ZN(n5514) );
  INVX0 U8053 ( .INP(n5515), .ZN(n5517) );
  INVX0 U8054 ( .INP(n5516), .ZN(n5518) );
  INVX0 U8055 ( .INP(n2912), .ZN(n5519) );
  INVX0 U8056 ( .INP(n5516), .ZN(n5520) );
  INVX0 U8057 ( .INP(n5527), .ZN(n5521) );
  INVX0 U8058 ( .INP(n2529), .ZN(n5528) );
  INVX0 U8059 ( .INP(n5536), .ZN(n5529) );
  INVX0 U8060 ( .INP(n5537), .ZN(n5530) );
  INVX0 U8061 ( .INP(n5535), .ZN(n5531) );
  INVX0 U8062 ( .INP(n5552), .ZN(n5539) );
  INVX0 U8063 ( .INP(n5552), .ZN(n5540) );
  INVX0 U8064 ( .INP(n5552), .ZN(n5541) );
  INVX0 U8065 ( .INP(n5552), .ZN(n5542) );
  INVX0 U8066 ( .INP(n5552), .ZN(n5543) );
  INVX0 U8067 ( .INP(n5552), .ZN(n5544) );
  NBUFFX2 U8068 ( .INP(n5550), .Z(n5545) );
  NBUFFX2 U8069 ( .INP(n5551), .Z(n5546) );
  NBUFFX2 U8070 ( .INP(n5550), .Z(n5547) );
  NBUFFX2 U8071 ( .INP(n5551), .Z(n5548) );
  NBUFFX2 U8072 ( .INP(n5550), .Z(n5549) );
  NBUFFX2 U8073 ( .INP(n4914), .Z(n5550) );
  NBUFFX2 U8074 ( .INP(n4914), .Z(n5551) );
  NBUFFX2 U8075 ( .INP(n4914), .Z(n5552) );
  INVX0 U8076 ( .INP(n5572), .ZN(n5553) );
  INVX0 U8077 ( .INP(n5562), .ZN(n5554) );
  INVX0 U8078 ( .INP(n5567), .ZN(n5555) );
  INVX0 U8079 ( .INP(n5566), .ZN(n5556) );
  INVX0 U8080 ( .INP(n5569), .ZN(n5557) );
  INVX0 U8081 ( .INP(n5564), .ZN(n5558) );
  INVX0 U8082 ( .INP(n5567), .ZN(n5559) );
  INVX0 U8083 ( .INP(n5564), .ZN(n5560) );
  INVX0 U8084 ( .INP(n5563), .ZN(n5561) );
  INVX0 U8085 ( .INP(n2525), .ZN(n5570) );
  INVX0 U8086 ( .INP(n2525), .ZN(n5571) );
  INVX0 U8087 ( .INP(n2525), .ZN(n5572) );
  INVX0 U8088 ( .INP(n5574), .ZN(n5576) );
  INVX0 U8089 ( .INP(n5575), .ZN(n5577) );
  INVX0 U8090 ( .INP(n2523), .ZN(n5578) );
  INVX0 U8091 ( .INP(n5585), .ZN(n5579) );
  INVX0 U8092 ( .INP(n5585), .ZN(n5580) );
  INVX0 U8093 ( .INP(n5591), .ZN(n5586) );
  INVX0 U8094 ( .INP(n5591), .ZN(n5587) );
  INVX0 U8095 ( .INP(n5591), .ZN(n5588) );
  INVX0 U8096 ( .INP(n5591), .ZN(n5589) );
  INVX0 U8097 ( .INP(n5591), .ZN(n5590) );
  INVX0 U8098 ( .INP(n1767), .ZN(n5600) );
  INVX0 U8099 ( .INP(n5610), .ZN(n5601) );
  INVX0 U8100 ( .INP(n5609), .ZN(n5602) );
  INVX0 U8101 ( .INP(n5597), .ZN(n5603) );
  INVX0 U8102 ( .INP(n5598), .ZN(n5604) );
  INVX0 U8103 ( .INP(n5598), .ZN(n5605) );
  INVX0 U8104 ( .INP(n5612), .ZN(n5606) );
  INVX0 U8105 ( .INP(n5599), .ZN(n5607) );
  INVX0 U8106 ( .INP(n5622), .ZN(n5616) );
  INVX0 U8107 ( .INP(n5622), .ZN(n5617) );
  INVX0 U8108 ( .INP(n5622), .ZN(n5618) );
  INVX0 U8109 ( .INP(n5622), .ZN(n5619) );
  INVX0 U8110 ( .INP(n5622), .ZN(n5620) );
  INVX0 U8111 ( .INP(n5622), .ZN(n5621) );
  INVX0 U8112 ( .INP(n1763), .ZN(n5624) );
  INVX0 U8113 ( .INP(n5636), .ZN(n5625) );
  INVX0 U8114 ( .INP(n5636), .ZN(n5626) );
  INVX0 U8115 ( .INP(n5636), .ZN(n5627) );
  INVX0 U8116 ( .INP(n5650), .ZN(n5637) );
  INVX0 U8117 ( .INP(n5648), .ZN(n5638) );
  INVX0 U8118 ( .INP(n4917), .ZN(n5639) );
  INVX0 U8119 ( .INP(n5647), .ZN(n5640) );
  INVX0 U8120 ( .INP(n5648), .ZN(n5641) );
  INVX0 U8121 ( .INP(n5644), .ZN(n5642) );
  NBUFFX2 U8122 ( .INP(n1759), .Z(n5651) );
  NBUFFX2 U8123 ( .INP(n1759), .Z(n5652) );
  INVX0 U8124 ( .INP(n5663), .ZN(n5653) );
  INVX0 U8125 ( .INP(n5663), .ZN(n5654) );
  INVX0 U8126 ( .INP(n5663), .ZN(n5655) );
  INVX0 U8127 ( .INP(n5663), .ZN(n5656) );
  INVX0 U8128 ( .INP(n5663), .ZN(n5657) );
  INVX0 U8129 ( .INP(n5663), .ZN(n5658) );
  INVX0 U8130 ( .INP(n5663), .ZN(n5659) );
  INVX0 U8131 ( .INP(n5663), .ZN(n5660) );
  INVX0 U8132 ( .INP(n5663), .ZN(n5661) );
  INVX0 U8133 ( .INP(n5663), .ZN(n5662) );
  NBUFFX2 U8134 ( .INP(n1759), .Z(n5663) );
  NBUFFX2 U8135 ( .INP(n5651), .Z(n5664) );
  NBUFFX2 U8136 ( .INP(n5651), .Z(n5665) );
  NBUFFX2 U8137 ( .INP(n5651), .Z(n5666) );
  NBUFFX2 U8138 ( .INP(n5651), .Z(n5667) );
  NBUFFX2 U8139 ( .INP(n5652), .Z(n5668) );
  NBUFFX2 U8140 ( .INP(n5652), .Z(n5669) );
  NBUFFX2 U8141 ( .INP(n5652), .Z(n5670) );
  INVX0 U8142 ( .INP(n5681), .ZN(n5671) );
  INVX0 U8143 ( .INP(n5677), .ZN(n5672) );
  INVX0 U8144 ( .INP(n1757), .ZN(n5673) );
  INVX0 U8145 ( .INP(n5676), .ZN(n5674) );
  INVX0 U8146 ( .INP(n5681), .ZN(n5675) );
  INVX0 U8147 ( .INP(n5684), .ZN(n5691) );
  INVX0 U8148 ( .INP(n5687), .ZN(n5692) );
  INVX0 U8149 ( .INP(n1124), .ZN(n5693) );
  INVX0 U8150 ( .INP(n5686), .ZN(n5694) );
  INVX0 U8151 ( .INP(n5688), .ZN(n5695) );
  INVX0 U8152 ( .INP(n5703), .ZN(n5696) );
  INVX0 U8153 ( .INP(n5707), .ZN(n5697) );
  INVX0 U8154 ( .INP(n5707), .ZN(n5698) );
  INVX0 U8155 ( .INP(n5707), .ZN(n5699) );
  INVX0 U8156 ( .INP(n5707), .ZN(n5700) );
  INVX0 U8157 ( .INP(n5707), .ZN(n5701) );
  NBUFFX2 U8158 ( .INP(n5201), .Z(n5702) );
  NBUFFX2 U8159 ( .INP(n5201), .Z(n5703) );
  NBUFFX2 U8160 ( .INP(n5201), .Z(n5704) );
  NBUFFX2 U8161 ( .INP(n5201), .Z(n5705) );
  NBUFFX2 U8162 ( .INP(n5201), .Z(n5706) );
  NBUFFX2 U8163 ( .INP(n5201), .Z(n5707) );
  INVX0 U8164 ( .INP(n4910), .ZN(n5708) );
  INVX0 U8165 ( .INP(n5719), .ZN(n5709) );
  INVX0 U8166 ( .INP(n5723), .ZN(n5710) );
  INVX0 U8167 ( .INP(n5726), .ZN(n5711) );
  INVX0 U8168 ( .INP(n5720), .ZN(n5712) );
  INVX0 U8169 ( .INP(n5719), .ZN(n5713) );
  INVX0 U8170 ( .INP(n5723), .ZN(n5714) );
  INVX0 U8171 ( .INP(n4910), .ZN(n5715) );
  INVX0 U8172 ( .INP(n5719), .ZN(n5716) );
  INVX0 U8173 ( .INP(n5740), .ZN(n5727) );
  INVX0 U8174 ( .INP(n5740), .ZN(n5728) );
  INVX0 U8175 ( .INP(n5740), .ZN(n5729) );
  INVX0 U8176 ( .INP(n5740), .ZN(n5730) );
  INVX0 U8177 ( .INP(n5740), .ZN(n5731) );
  INVX0 U8178 ( .INP(n5740), .ZN(n5732) );
  NBUFFX2 U8179 ( .INP(n5738), .Z(n5733) );
  NBUFFX2 U8180 ( .INP(n5739), .Z(n5734) );
  NBUFFX2 U8181 ( .INP(n5738), .Z(n5735) );
  NBUFFX2 U8182 ( .INP(n5739), .Z(n5736) );
  NBUFFX2 U8183 ( .INP(n5738), .Z(n5737) );
  NBUFFX2 U8184 ( .INP(n4915), .Z(n5738) );
  NBUFFX2 U8185 ( .INP(n4915), .Z(n5739) );
  NBUFFX2 U8186 ( .INP(n4915), .Z(n5740) );
  INVX0 U8187 ( .INP(n5760), .ZN(n5741) );
  INVX0 U8188 ( .INP(n5750), .ZN(n5742) );
  INVX0 U8189 ( .INP(n5755), .ZN(n5743) );
  INVX0 U8190 ( .INP(n5754), .ZN(n5744) );
  INVX0 U8191 ( .INP(n5757), .ZN(n5745) );
  INVX0 U8192 ( .INP(n5752), .ZN(n5746) );
  INVX0 U8193 ( .INP(n5755), .ZN(n5747) );
  INVX0 U8194 ( .INP(n5752), .ZN(n5748) );
  INVX0 U8195 ( .INP(n5751), .ZN(n5749) );
  INVX0 U8196 ( .INP(n1116), .ZN(n5758) );
  INVX0 U8197 ( .INP(n1116), .ZN(n5759) );
  INVX0 U8198 ( .INP(n1116), .ZN(n5760) );
  INVX0 U8199 ( .INP(n5766), .ZN(n5761) );
  INVX0 U8200 ( .INP(n5766), .ZN(n5762) );
  INVX0 U8201 ( .INP(n5766), .ZN(n5763) );
  INVX0 U8202 ( .INP(n5766), .ZN(n5764) );
  INVX0 U8203 ( .INP(n5766), .ZN(n5765) );
  INVX0 U8204 ( .INP(n5783), .ZN(n5773) );
  INVX0 U8205 ( .INP(n5781), .ZN(n5774) );
  INVX0 U8206 ( .INP(n5785), .ZN(n5775) );
  INVX0 U8207 ( .INP(n5786), .ZN(n5776) );
  INVX0 U8208 ( .INP(n5784), .ZN(n5777) );
  INVX0 U8209 ( .INP(n4919), .ZN(n5778) );
  INVX0 U8210 ( .INP(n5789), .ZN(n5790) );
  INVX0 U8211 ( .INP(n5788), .ZN(n5791) );
  INVX0 U8212 ( .INP(n5787), .ZN(n5792) );
  INVX0 U8213 ( .INP(n5807), .ZN(n5793) );
  INVX0 U8214 ( .INP(n5806), .ZN(n5794) );
  INVX0 U8215 ( .INP(n5789), .ZN(n5795) );
  INVX0 U8216 ( .INP(n5787), .ZN(n5796) );
  INVX0 U8217 ( .INP(n5789), .ZN(n5797) );
  INVX0 U8218 ( .INP(n5802), .ZN(n5798) );
  INVX0 U8219 ( .INP(n5800), .ZN(n5799) );
  INVX0 U8220 ( .INP(n5817), .ZN(n5808) );
  INVX0 U8221 ( .INP(n5821), .ZN(n5809) );
  INVX0 U8222 ( .INP(n4918), .ZN(n5810) );
  INVX0 U8223 ( .INP(n5814), .ZN(n5811) );
  INVX0 U8224 ( .INP(n5821), .ZN(n5812) );
  INVX0 U8225 ( .INP(n5818), .ZN(n5813) );
  INVX0 U8226 ( .INP(n5825), .ZN(n5826) );
  INVX0 U8227 ( .INP(n5836), .ZN(n5827) );
  INVX0 U8228 ( .INP(n5824), .ZN(n5828) );
  INVX0 U8229 ( .INP(n5822), .ZN(n5829) );
  INVX0 U8230 ( .INP(n5842), .ZN(n5830) );
  INVX0 U8231 ( .INP(n5838), .ZN(n5831) );
  INVX0 U8232 ( .INP(n5824), .ZN(n5832) );
  INVX0 U8233 ( .INP(n5841), .ZN(n5833) );
  INVX0 U8234 ( .INP(n5837), .ZN(n5834) );
  INVX0 U8235 ( .INP(n5840), .ZN(n5835) );
  INVX0 U8236 ( .INP(n5852), .ZN(n5843) );
  INVX0 U8237 ( .INP(n5851), .ZN(n5844) );
  INVX0 U8238 ( .INP(n826), .ZN(n5845) );
  INVX0 U8239 ( .INP(n5852), .ZN(n5846) );
  INVX0 U8240 ( .INP(n5849), .ZN(n5847) );
  INVX0 U8241 ( .INP(\decodedPacket[2][121] ), .ZN(n5854) );
  INVX0 U8242 ( .INP(\decodedPacket[6][121] ), .ZN(n5856) );
  XOR2X1 U8243 ( .IN1(\add_177_I7_aco/carry[5] ), .IN2(N6449), .Q(N8585) );
  AND2X1 U8244 ( .IN1(N6448), .IN2(\add_177_I7_aco/carry[4] ), .Q(
        \add_177_I7_aco/carry[5] ) );
  XOR2X1 U8245 ( .IN1(\add_177_I7_aco/carry[4] ), .IN2(N6448), .Q(N8584) );
  AND2X1 U8246 ( .IN1(N6447), .IN2(\add_177_I7_aco/carry[3] ), .Q(
        \add_177_I7_aco/carry[4] ) );
  XOR2X1 U8247 ( .IN1(\add_177_I7_aco/carry[3] ), .IN2(N6447), .Q(N8583) );
  AND2X1 U8248 ( .IN1(N6446), .IN2(\add_177_I7_aco/carry[2] ), .Q(
        \add_177_I7_aco/carry[3] ) );
  XOR2X1 U8249 ( .IN1(\add_177_I7_aco/carry[2] ), .IN2(N6446), .Q(N8582) );
  AND2X1 U8250 ( .IN1(N6445), .IN2(\add_177_I7_aco/carry[1] ), .Q(
        \add_177_I7_aco/carry[2] ) );
  XOR2X1 U8251 ( .IN1(\add_177_I7_aco/carry[1] ), .IN2(N6445), .Q(N8581) );
  AND2X1 U8252 ( .IN1(N6444), .IN2(decodedPacketValid[6]), .Q(
        \add_177_I7_aco/carry[1] ) );
  XOR2X1 U8253 ( .IN1(decodedPacketValid[6]), .IN2(N6444), .Q(N8580) );
  AND2X1 U8254 ( .IN1(N4312), .IN2(\add_177_I6_aco/carry[4] ), .Q(N6449) );
  XOR2X1 U8255 ( .IN1(\add_177_I6_aco/carry[4] ), .IN2(N4312), .Q(N6448) );
  AND2X1 U8256 ( .IN1(N4311), .IN2(\add_177_I6_aco/carry[3] ), .Q(
        \add_177_I6_aco/carry[4] ) );
  XOR2X1 U8257 ( .IN1(\add_177_I6_aco/carry[3] ), .IN2(N4311), .Q(N6447) );
  AND2X1 U8258 ( .IN1(N2175), .IN2(\add_177_I5_aco/carry[3] ), .Q(N4312) );
  XOR2X1 U8259 ( .IN1(\add_177_I5_aco/carry[3] ), .IN2(N2175), .Q(N4311) );
  AND2X1 U8260 ( .IN1(N4310), .IN2(\add_177_I6_aco/carry[2] ), .Q(
        \add_177_I6_aco/carry[3] ) );
  XOR2X1 U8261 ( .IN1(\add_177_I6_aco/carry[2] ), .IN2(N4310), .Q(N6446) );
  AND2X1 U8262 ( .IN1(N2174), .IN2(\add_177_I5_aco/carry[2] ), .Q(
        \add_177_I5_aco/carry[3] ) );
  XOR2X1 U8263 ( .IN1(\add_177_I5_aco/carry[2] ), .IN2(N2174), .Q(N4310) );
  AND2X1 U8264 ( .IN1(N1070), .IN2(\add_177_I4_aco/carry[2] ), .Q(N2175) );
  XOR2X1 U8265 ( .IN1(\add_177_I4_aco/carry[2] ), .IN2(N1070), .Q(N2174) );
  AND2X1 U8266 ( .IN1(N4309), .IN2(\add_177_I6_aco/carry[1] ), .Q(
        \add_177_I6_aco/carry[2] ) );
  XOR2X1 U8267 ( .IN1(\add_177_I6_aco/carry[1] ), .IN2(N4309), .Q(N6445) );
  AND2X1 U8268 ( .IN1(N4308), .IN2(decodedPacketValid[5]), .Q(
        \add_177_I6_aco/carry[1] ) );
  XOR2X1 U8269 ( .IN1(decodedPacketValid[5]), .IN2(N4308), .Q(N6444) );
  AND2X1 U8270 ( .IN1(N2173), .IN2(\add_177_I5_aco/carry[1] ), .Q(
        \add_177_I5_aco/carry[2] ) );
  XOR2X1 U8271 ( .IN1(\add_177_I5_aco/carry[1] ), .IN2(N2173), .Q(N4309) );
  AND2X1 U8272 ( .IN1(N2172), .IN2(decodedPacketValid[4]), .Q(
        \add_177_I5_aco/carry[1] ) );
  XOR2X1 U8273 ( .IN1(decodedPacketValid[4]), .IN2(N2172), .Q(N4308) );
  AND2X1 U8274 ( .IN1(N1069), .IN2(\add_177_I4_aco/carry[1] ), .Q(
        \add_177_I4_aco/carry[2] ) );
  XOR2X1 U8275 ( .IN1(\add_177_I4_aco/carry[1] ), .IN2(N1069), .Q(N2173) );
  AND2X1 U8276 ( .IN1(N1068), .IN2(decodedPacketValid[3]), .Q(
        \add_177_I4_aco/carry[1] ) );
  XOR2X1 U8277 ( .IN1(decodedPacketValid[3]), .IN2(N1068), .Q(N2172) );
  AND2X1 U8278 ( .IN1(\add_177_I3_aco/A[1] ), .IN2(\add_177_I3_aco/carry[1] ), 
        .Q(N1070) );
  XOR2X1 U8279 ( .IN1(\add_177_I3_aco/carry[1] ), .IN2(\add_177_I3_aco/A[1] ), 
        .Q(N1069) );
  AND2X1 U8280 ( .IN1(\add_177_I3_aco/A[0] ), .IN2(decodedPacketValid[2]), .Q(
        \add_177_I3_aco/carry[1] ) );
  XOR2X1 U8281 ( .IN1(decodedPacketValid[2]), .IN2(\add_177_I3_aco/A[0] ), .Q(
        N1068) );
endmodule

